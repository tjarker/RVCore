module IF(
  input         clock,
  input         reset,
  input  [31:0] in_pcNext,
  input         in_branch,
  output [31:0] out_pc,
  output [31:0] out_instr,
  input         ctrl_pcEn
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[IF.scala 18:19]
  wire [31:0] _T_1 = pc + 32'h3; // @[IF.scala 28:27]
  wire [31:0] _T_4 = pc + 32'h2; // @[IF.scala 28:43]
  wire [31:0] _T_7 = pc + 32'h1; // @[IF.scala 28:59]
  wire [7:0] _GEN_1 = 10'h1 == _T_7[9:0] ? 8'h21 : 8'h97; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2 = 10'h2 == _T_7[9:0] ? 8'h0 : _GEN_1; // @[Cat.scala 29:58]
  wire [7:0] _GEN_3 = 10'h3 == _T_7[9:0] ? 8'h0 : _GEN_2; // @[Cat.scala 29:58]
  wire [7:0] _GEN_4 = 10'h4 == _T_7[9:0] ? 8'h93 : _GEN_3; // @[Cat.scala 29:58]
  wire [7:0] _GEN_5 = 10'h5 == _T_7[9:0] ? 8'h81 : _GEN_4; // @[Cat.scala 29:58]
  wire [7:0] _GEN_6 = 10'h6 == _T_7[9:0] ? 8'h1 : _GEN_5; // @[Cat.scala 29:58]
  wire [7:0] _GEN_7 = 10'h7 == _T_7[9:0] ? 8'h97 : _GEN_6; // @[Cat.scala 29:58]
  wire [7:0] _GEN_8 = 10'h8 == _T_7[9:0] ? 8'h17 : _GEN_7; // @[Cat.scala 29:58]
  wire [7:0] _GEN_9 = 10'h9 == _T_7[9:0] ? 8'h11 : _GEN_8; // @[Cat.scala 29:58]
  wire [7:0] _GEN_10 = 10'ha == _T_7[9:0] ? 8'h0 : _GEN_9; // @[Cat.scala 29:58]
  wire [7:0] _GEN_11 = 10'hb == _T_7[9:0] ? 8'h0 : _GEN_10; // @[Cat.scala 29:58]
  wire [7:0] _GEN_12 = 10'hc == _T_7[9:0] ? 8'h13 : _GEN_11; // @[Cat.scala 29:58]
  wire [7:0] _GEN_13 = 10'hd == _T_7[9:0] ? 8'h1 : _GEN_12; // @[Cat.scala 29:58]
  wire [7:0] _GEN_14 = 10'he == _T_7[9:0] ? 8'h81 : _GEN_13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_15 = 10'hf == _T_7[9:0] ? 8'hff : _GEN_14; // @[Cat.scala 29:58]
  wire [7:0] _GEN_16 = 10'h10 == _T_7[9:0] ? 8'h33 : _GEN_15; // @[Cat.scala 29:58]
  wire [7:0] _GEN_17 = 10'h11 == _T_7[9:0] ? 8'h4 : _GEN_16; // @[Cat.scala 29:58]
  wire [7:0] _GEN_18 = 10'h12 == _T_7[9:0] ? 8'h1 : _GEN_17; // @[Cat.scala 29:58]
  wire [7:0] _GEN_19 = 10'h13 == _T_7[9:0] ? 8'h0 : _GEN_18; // @[Cat.scala 29:58]
  wire [7:0] _GEN_20 = 10'h14 == _T_7[9:0] ? 8'h6f : _GEN_19; // @[Cat.scala 29:58]
  wire [7:0] _GEN_21 = 10'h15 == _T_7[9:0] ? 8'h0 : _GEN_20; // @[Cat.scala 29:58]
  wire [7:0] _GEN_22 = 10'h16 == _T_7[9:0] ? 8'h80 : _GEN_21; // @[Cat.scala 29:58]
  wire [7:0] _GEN_23 = 10'h17 == _T_7[9:0] ? 8'h9 : _GEN_22; // @[Cat.scala 29:58]
  wire [7:0] _GEN_24 = 10'h18 == _T_7[9:0] ? 8'h13 : _GEN_23; // @[Cat.scala 29:58]
  wire [7:0] _GEN_25 = 10'h19 == _T_7[9:0] ? 8'h1 : _GEN_24; // @[Cat.scala 29:58]
  wire [7:0] _GEN_26 = 10'h1a == _T_7[9:0] ? 8'h1 : _GEN_25; // @[Cat.scala 29:58]
  wire [7:0] _GEN_27 = 10'h1b == _T_7[9:0] ? 8'hfe : _GEN_26; // @[Cat.scala 29:58]
  wire [7:0] _GEN_28 = 10'h1c == _T_7[9:0] ? 8'h23 : _GEN_27; // @[Cat.scala 29:58]
  wire [7:0] _GEN_29 = 10'h1d == _T_7[9:0] ? 8'h2e : _GEN_28; // @[Cat.scala 29:58]
  wire [7:0] _GEN_30 = 10'h1e == _T_7[9:0] ? 8'h81 : _GEN_29; // @[Cat.scala 29:58]
  wire [7:0] _GEN_31 = 10'h1f == _T_7[9:0] ? 8'h0 : _GEN_30; // @[Cat.scala 29:58]
  wire [7:0] _GEN_32 = 10'h20 == _T_7[9:0] ? 8'h13 : _GEN_31; // @[Cat.scala 29:58]
  wire [7:0] _GEN_33 = 10'h21 == _T_7[9:0] ? 8'h4 : _GEN_32; // @[Cat.scala 29:58]
  wire [7:0] _GEN_34 = 10'h22 == _T_7[9:0] ? 8'h1 : _GEN_33; // @[Cat.scala 29:58]
  wire [7:0] _GEN_35 = 10'h23 == _T_7[9:0] ? 8'h2 : _GEN_34; // @[Cat.scala 29:58]
  wire [7:0] _GEN_36 = 10'h24 == _T_7[9:0] ? 8'hb7 : _GEN_35; // @[Cat.scala 29:58]
  wire [7:0] _GEN_37 = 10'h25 == _T_7[9:0] ? 8'h27 : _GEN_36; // @[Cat.scala 29:58]
  wire [7:0] _GEN_38 = 10'h26 == _T_7[9:0] ? 8'h0 : _GEN_37; // @[Cat.scala 29:58]
  wire [7:0] _GEN_39 = 10'h27 == _T_7[9:0] ? 8'h0 : _GEN_38; // @[Cat.scala 29:58]
  wire [7:0] _GEN_40 = 10'h28 == _T_7[9:0] ? 8'h93 : _GEN_39; // @[Cat.scala 29:58]
  wire [7:0] _GEN_41 = 10'h29 == _T_7[9:0] ? 8'h87 : _GEN_40; // @[Cat.scala 29:58]
  wire [7:0] _GEN_42 = 10'h2a == _T_7[9:0] ? 8'h7 : _GEN_41; // @[Cat.scala 29:58]
  wire [7:0] _GEN_43 = 10'h2b == _T_7[9:0] ? 8'h20 : _GEN_42; // @[Cat.scala 29:58]
  wire [7:0] _GEN_44 = 10'h2c == _T_7[9:0] ? 8'h23 : _GEN_43; // @[Cat.scala 29:58]
  wire [7:0] _GEN_45 = 10'h2d == _T_7[9:0] ? 8'h26 : _GEN_44; // @[Cat.scala 29:58]
  wire [7:0] _GEN_46 = 10'h2e == _T_7[9:0] ? 8'hf4 : _GEN_45; // @[Cat.scala 29:58]
  wire [7:0] _GEN_47 = 10'h2f == _T_7[9:0] ? 8'hfe : _GEN_46; // @[Cat.scala 29:58]
  wire [7:0] _GEN_48 = 10'h30 == _T_7[9:0] ? 8'h83 : _GEN_47; // @[Cat.scala 29:58]
  wire [7:0] _GEN_49 = 10'h31 == _T_7[9:0] ? 8'h27 : _GEN_48; // @[Cat.scala 29:58]
  wire [7:0] _GEN_50 = 10'h32 == _T_7[9:0] ? 8'hc4 : _GEN_49; // @[Cat.scala 29:58]
  wire [7:0] _GEN_51 = 10'h33 == _T_7[9:0] ? 8'hfe : _GEN_50; // @[Cat.scala 29:58]
  wire [7:0] _GEN_52 = 10'h34 == _T_7[9:0] ? 8'h83 : _GEN_51; // @[Cat.scala 29:58]
  wire [7:0] _GEN_53 = 10'h35 == _T_7[9:0] ? 8'ha7 : _GEN_52; // @[Cat.scala 29:58]
  wire [7:0] _GEN_54 = 10'h36 == _T_7[9:0] ? 8'h7 : _GEN_53; // @[Cat.scala 29:58]
  wire [7:0] _GEN_55 = 10'h37 == _T_7[9:0] ? 8'h0 : _GEN_54; // @[Cat.scala 29:58]
  wire [7:0] _GEN_56 = 10'h38 == _T_7[9:0] ? 8'h13 : _GEN_55; // @[Cat.scala 29:58]
  wire [7:0] _GEN_57 = 10'h39 == _T_7[9:0] ? 8'h85 : _GEN_56; // @[Cat.scala 29:58]
  wire [7:0] _GEN_58 = 10'h3a == _T_7[9:0] ? 8'h7 : _GEN_57; // @[Cat.scala 29:58]
  wire [7:0] _GEN_59 = 10'h3b == _T_7[9:0] ? 8'h0 : _GEN_58; // @[Cat.scala 29:58]
  wire [7:0] _GEN_60 = 10'h3c == _T_7[9:0] ? 8'h3 : _GEN_59; // @[Cat.scala 29:58]
  wire [7:0] _GEN_61 = 10'h3d == _T_7[9:0] ? 8'h24 : _GEN_60; // @[Cat.scala 29:58]
  wire [7:0] _GEN_62 = 10'h3e == _T_7[9:0] ? 8'hc1 : _GEN_61; // @[Cat.scala 29:58]
  wire [7:0] _GEN_63 = 10'h3f == _T_7[9:0] ? 8'h1 : _GEN_62; // @[Cat.scala 29:58]
  wire [7:0] _GEN_64 = 10'h40 == _T_7[9:0] ? 8'h13 : _GEN_63; // @[Cat.scala 29:58]
  wire [7:0] _GEN_65 = 10'h41 == _T_7[9:0] ? 8'h1 : _GEN_64; // @[Cat.scala 29:58]
  wire [7:0] _GEN_66 = 10'h42 == _T_7[9:0] ? 8'h1 : _GEN_65; // @[Cat.scala 29:58]
  wire [7:0] _GEN_67 = 10'h43 == _T_7[9:0] ? 8'h2 : _GEN_66; // @[Cat.scala 29:58]
  wire [7:0] _GEN_68 = 10'h44 == _T_7[9:0] ? 8'h67 : _GEN_67; // @[Cat.scala 29:58]
  wire [7:0] _GEN_69 = 10'h45 == _T_7[9:0] ? 8'h80 : _GEN_68; // @[Cat.scala 29:58]
  wire [7:0] _GEN_70 = 10'h46 == _T_7[9:0] ? 8'h0 : _GEN_69; // @[Cat.scala 29:58]
  wire [7:0] _GEN_71 = 10'h47 == _T_7[9:0] ? 8'h0 : _GEN_70; // @[Cat.scala 29:58]
  wire [7:0] _GEN_72 = 10'h48 == _T_7[9:0] ? 8'h13 : _GEN_71; // @[Cat.scala 29:58]
  wire [7:0] _GEN_73 = 10'h49 == _T_7[9:0] ? 8'h1 : _GEN_72; // @[Cat.scala 29:58]
  wire [7:0] _GEN_74 = 10'h4a == _T_7[9:0] ? 8'h1 : _GEN_73; // @[Cat.scala 29:58]
  wire [7:0] _GEN_75 = 10'h4b == _T_7[9:0] ? 8'hfe : _GEN_74; // @[Cat.scala 29:58]
  wire [7:0] _GEN_76 = 10'h4c == _T_7[9:0] ? 8'h23 : _GEN_75; // @[Cat.scala 29:58]
  wire [7:0] _GEN_77 = 10'h4d == _T_7[9:0] ? 8'h2e : _GEN_76; // @[Cat.scala 29:58]
  wire [7:0] _GEN_78 = 10'h4e == _T_7[9:0] ? 8'h81 : _GEN_77; // @[Cat.scala 29:58]
  wire [7:0] _GEN_79 = 10'h4f == _T_7[9:0] ? 8'h0 : _GEN_78; // @[Cat.scala 29:58]
  wire [7:0] _GEN_80 = 10'h50 == _T_7[9:0] ? 8'h13 : _GEN_79; // @[Cat.scala 29:58]
  wire [7:0] _GEN_81 = 10'h51 == _T_7[9:0] ? 8'h4 : _GEN_80; // @[Cat.scala 29:58]
  wire [7:0] _GEN_82 = 10'h52 == _T_7[9:0] ? 8'h1 : _GEN_81; // @[Cat.scala 29:58]
  wire [7:0] _GEN_83 = 10'h53 == _T_7[9:0] ? 8'h2 : _GEN_82; // @[Cat.scala 29:58]
  wire [7:0] _GEN_84 = 10'h54 == _T_7[9:0] ? 8'hb7 : _GEN_83; // @[Cat.scala 29:58]
  wire [7:0] _GEN_85 = 10'h55 == _T_7[9:0] ? 8'h27 : _GEN_84; // @[Cat.scala 29:58]
  wire [7:0] _GEN_86 = 10'h56 == _T_7[9:0] ? 8'h0 : _GEN_85; // @[Cat.scala 29:58]
  wire [7:0] _GEN_87 = 10'h57 == _T_7[9:0] ? 8'h0 : _GEN_86; // @[Cat.scala 29:58]
  wire [7:0] _GEN_88 = 10'h58 == _T_7[9:0] ? 8'h93 : _GEN_87; // @[Cat.scala 29:58]
  wire [7:0] _GEN_89 = 10'h59 == _T_7[9:0] ? 8'h87 : _GEN_88; // @[Cat.scala 29:58]
  wire [7:0] _GEN_90 = 10'h5a == _T_7[9:0] ? 8'h7 : _GEN_89; // @[Cat.scala 29:58]
  wire [7:0] _GEN_91 = 10'h5b == _T_7[9:0] ? 8'h10 : _GEN_90; // @[Cat.scala 29:58]
  wire [7:0] _GEN_92 = 10'h5c == _T_7[9:0] ? 8'h23 : _GEN_91; // @[Cat.scala 29:58]
  wire [7:0] _GEN_93 = 10'h5d == _T_7[9:0] ? 8'h26 : _GEN_92; // @[Cat.scala 29:58]
  wire [7:0] _GEN_94 = 10'h5e == _T_7[9:0] ? 8'hf4 : _GEN_93; // @[Cat.scala 29:58]
  wire [7:0] _GEN_95 = 10'h5f == _T_7[9:0] ? 8'hfe : _GEN_94; // @[Cat.scala 29:58]
  wire [7:0] _GEN_96 = 10'h60 == _T_7[9:0] ? 8'h83 : _GEN_95; // @[Cat.scala 29:58]
  wire [7:0] _GEN_97 = 10'h61 == _T_7[9:0] ? 8'h27 : _GEN_96; // @[Cat.scala 29:58]
  wire [7:0] _GEN_98 = 10'h62 == _T_7[9:0] ? 8'hc4 : _GEN_97; // @[Cat.scala 29:58]
  wire [7:0] _GEN_99 = 10'h63 == _T_7[9:0] ? 8'hfe : _GEN_98; // @[Cat.scala 29:58]
  wire [7:0] _GEN_100 = 10'h64 == _T_7[9:0] ? 8'h83 : _GEN_99; // @[Cat.scala 29:58]
  wire [7:0] _GEN_101 = 10'h65 == _T_7[9:0] ? 8'ha7 : _GEN_100; // @[Cat.scala 29:58]
  wire [7:0] _GEN_102 = 10'h66 == _T_7[9:0] ? 8'h7 : _GEN_101; // @[Cat.scala 29:58]
  wire [7:0] _GEN_103 = 10'h67 == _T_7[9:0] ? 8'h0 : _GEN_102; // @[Cat.scala 29:58]
  wire [7:0] _GEN_104 = 10'h68 == _T_7[9:0] ? 8'h13 : _GEN_103; // @[Cat.scala 29:58]
  wire [7:0] _GEN_105 = 10'h69 == _T_7[9:0] ? 8'h85 : _GEN_104; // @[Cat.scala 29:58]
  wire [7:0] _GEN_106 = 10'h6a == _T_7[9:0] ? 8'h7 : _GEN_105; // @[Cat.scala 29:58]
  wire [7:0] _GEN_107 = 10'h6b == _T_7[9:0] ? 8'h0 : _GEN_106; // @[Cat.scala 29:58]
  wire [7:0] _GEN_108 = 10'h6c == _T_7[9:0] ? 8'h3 : _GEN_107; // @[Cat.scala 29:58]
  wire [7:0] _GEN_109 = 10'h6d == _T_7[9:0] ? 8'h24 : _GEN_108; // @[Cat.scala 29:58]
  wire [7:0] _GEN_110 = 10'h6e == _T_7[9:0] ? 8'hc1 : _GEN_109; // @[Cat.scala 29:58]
  wire [7:0] _GEN_111 = 10'h6f == _T_7[9:0] ? 8'h1 : _GEN_110; // @[Cat.scala 29:58]
  wire [7:0] _GEN_112 = 10'h70 == _T_7[9:0] ? 8'h13 : _GEN_111; // @[Cat.scala 29:58]
  wire [7:0] _GEN_113 = 10'h71 == _T_7[9:0] ? 8'h1 : _GEN_112; // @[Cat.scala 29:58]
  wire [7:0] _GEN_114 = 10'h72 == _T_7[9:0] ? 8'h1 : _GEN_113; // @[Cat.scala 29:58]
  wire [7:0] _GEN_115 = 10'h73 == _T_7[9:0] ? 8'h2 : _GEN_114; // @[Cat.scala 29:58]
  wire [7:0] _GEN_116 = 10'h74 == _T_7[9:0] ? 8'h67 : _GEN_115; // @[Cat.scala 29:58]
  wire [7:0] _GEN_117 = 10'h75 == _T_7[9:0] ? 8'h80 : _GEN_116; // @[Cat.scala 29:58]
  wire [7:0] _GEN_118 = 10'h76 == _T_7[9:0] ? 8'h0 : _GEN_117; // @[Cat.scala 29:58]
  wire [7:0] _GEN_119 = 10'h77 == _T_7[9:0] ? 8'h0 : _GEN_118; // @[Cat.scala 29:58]
  wire [7:0] _GEN_120 = 10'h78 == _T_7[9:0] ? 8'h13 : _GEN_119; // @[Cat.scala 29:58]
  wire [7:0] _GEN_121 = 10'h79 == _T_7[9:0] ? 8'h1 : _GEN_120; // @[Cat.scala 29:58]
  wire [7:0] _GEN_122 = 10'h7a == _T_7[9:0] ? 8'h1 : _GEN_121; // @[Cat.scala 29:58]
  wire [7:0] _GEN_123 = 10'h7b == _T_7[9:0] ? 8'hfd : _GEN_122; // @[Cat.scala 29:58]
  wire [7:0] _GEN_124 = 10'h7c == _T_7[9:0] ? 8'h23 : _GEN_123; // @[Cat.scala 29:58]
  wire [7:0] _GEN_125 = 10'h7d == _T_7[9:0] ? 8'h26 : _GEN_124; // @[Cat.scala 29:58]
  wire [7:0] _GEN_126 = 10'h7e == _T_7[9:0] ? 8'h81 : _GEN_125; // @[Cat.scala 29:58]
  wire [7:0] _GEN_127 = 10'h7f == _T_7[9:0] ? 8'h2 : _GEN_126; // @[Cat.scala 29:58]
  wire [7:0] _GEN_128 = 10'h80 == _T_7[9:0] ? 8'h13 : _GEN_127; // @[Cat.scala 29:58]
  wire [7:0] _GEN_129 = 10'h81 == _T_7[9:0] ? 8'h4 : _GEN_128; // @[Cat.scala 29:58]
  wire [7:0] _GEN_130 = 10'h82 == _T_7[9:0] ? 8'h1 : _GEN_129; // @[Cat.scala 29:58]
  wire [7:0] _GEN_131 = 10'h83 == _T_7[9:0] ? 8'h3 : _GEN_130; // @[Cat.scala 29:58]
  wire [7:0] _GEN_132 = 10'h84 == _T_7[9:0] ? 8'h23 : _GEN_131; // @[Cat.scala 29:58]
  wire [7:0] _GEN_133 = 10'h85 == _T_7[9:0] ? 8'h2e : _GEN_132; // @[Cat.scala 29:58]
  wire [7:0] _GEN_134 = 10'h86 == _T_7[9:0] ? 8'ha4 : _GEN_133; // @[Cat.scala 29:58]
  wire [7:0] _GEN_135 = 10'h87 == _T_7[9:0] ? 8'hfc : _GEN_134; // @[Cat.scala 29:58]
  wire [7:0] _GEN_136 = 10'h88 == _T_7[9:0] ? 8'hb7 : _GEN_135; // @[Cat.scala 29:58]
  wire [7:0] _GEN_137 = 10'h89 == _T_7[9:0] ? 8'h27 : _GEN_136; // @[Cat.scala 29:58]
  wire [7:0] _GEN_138 = 10'h8a == _T_7[9:0] ? 8'h0 : _GEN_137; // @[Cat.scala 29:58]
  wire [7:0] _GEN_139 = 10'h8b == _T_7[9:0] ? 8'h0 : _GEN_138; // @[Cat.scala 29:58]
  wire [7:0] _GEN_140 = 10'h8c == _T_7[9:0] ? 8'h23 : _GEN_139; // @[Cat.scala 29:58]
  wire [7:0] _GEN_141 = 10'h8d == _T_7[9:0] ? 8'h26 : _GEN_140; // @[Cat.scala 29:58]
  wire [7:0] _GEN_142 = 10'h8e == _T_7[9:0] ? 8'hf4 : _GEN_141; // @[Cat.scala 29:58]
  wire [7:0] _GEN_143 = 10'h8f == _T_7[9:0] ? 8'hfe : _GEN_142; // @[Cat.scala 29:58]
  wire [7:0] _GEN_144 = 10'h90 == _T_7[9:0] ? 8'h83 : _GEN_143; // @[Cat.scala 29:58]
  wire [7:0] _GEN_145 = 10'h91 == _T_7[9:0] ? 8'h27 : _GEN_144; // @[Cat.scala 29:58]
  wire [7:0] _GEN_146 = 10'h92 == _T_7[9:0] ? 8'hc4 : _GEN_145; // @[Cat.scala 29:58]
  wire [7:0] _GEN_147 = 10'h93 == _T_7[9:0] ? 8'hfe : _GEN_146; // @[Cat.scala 29:58]
  wire [7:0] _GEN_148 = 10'h94 == _T_7[9:0] ? 8'h3 : _GEN_147; // @[Cat.scala 29:58]
  wire [7:0] _GEN_149 = 10'h95 == _T_7[9:0] ? 8'h27 : _GEN_148; // @[Cat.scala 29:58]
  wire [7:0] _GEN_150 = 10'h96 == _T_7[9:0] ? 8'hc4 : _GEN_149; // @[Cat.scala 29:58]
  wire [7:0] _GEN_151 = 10'h97 == _T_7[9:0] ? 8'hfd : _GEN_150; // @[Cat.scala 29:58]
  wire [7:0] _GEN_152 = 10'h98 == _T_7[9:0] ? 8'h23 : _GEN_151; // @[Cat.scala 29:58]
  wire [7:0] _GEN_153 = 10'h99 == _T_7[9:0] ? 8'ha0 : _GEN_152; // @[Cat.scala 29:58]
  wire [7:0] _GEN_154 = 10'h9a == _T_7[9:0] ? 8'he7 : _GEN_153; // @[Cat.scala 29:58]
  wire [7:0] _GEN_155 = 10'h9b == _T_7[9:0] ? 8'h0 : _GEN_154; // @[Cat.scala 29:58]
  wire [7:0] _GEN_156 = 10'h9c == _T_7[9:0] ? 8'h13 : _GEN_155; // @[Cat.scala 29:58]
  wire [7:0] _GEN_157 = 10'h9d == _T_7[9:0] ? 8'h0 : _GEN_156; // @[Cat.scala 29:58]
  wire [7:0] _GEN_158 = 10'h9e == _T_7[9:0] ? 8'h0 : _GEN_157; // @[Cat.scala 29:58]
  wire [7:0] _GEN_159 = 10'h9f == _T_7[9:0] ? 8'h0 : _GEN_158; // @[Cat.scala 29:58]
  wire [7:0] _GEN_160 = 10'ha0 == _T_7[9:0] ? 8'h3 : _GEN_159; // @[Cat.scala 29:58]
  wire [7:0] _GEN_161 = 10'ha1 == _T_7[9:0] ? 8'h24 : _GEN_160; // @[Cat.scala 29:58]
  wire [7:0] _GEN_162 = 10'ha2 == _T_7[9:0] ? 8'hc1 : _GEN_161; // @[Cat.scala 29:58]
  wire [7:0] _GEN_163 = 10'ha3 == _T_7[9:0] ? 8'h2 : _GEN_162; // @[Cat.scala 29:58]
  wire [7:0] _GEN_164 = 10'ha4 == _T_7[9:0] ? 8'h13 : _GEN_163; // @[Cat.scala 29:58]
  wire [7:0] _GEN_165 = 10'ha5 == _T_7[9:0] ? 8'h1 : _GEN_164; // @[Cat.scala 29:58]
  wire [7:0] _GEN_166 = 10'ha6 == _T_7[9:0] ? 8'h1 : _GEN_165; // @[Cat.scala 29:58]
  wire [7:0] _GEN_167 = 10'ha7 == _T_7[9:0] ? 8'h3 : _GEN_166; // @[Cat.scala 29:58]
  wire [7:0] _GEN_168 = 10'ha8 == _T_7[9:0] ? 8'h67 : _GEN_167; // @[Cat.scala 29:58]
  wire [7:0] _GEN_169 = 10'ha9 == _T_7[9:0] ? 8'h80 : _GEN_168; // @[Cat.scala 29:58]
  wire [7:0] _GEN_170 = 10'haa == _T_7[9:0] ? 8'h0 : _GEN_169; // @[Cat.scala 29:58]
  wire [7:0] _GEN_171 = 10'hab == _T_7[9:0] ? 8'h0 : _GEN_170; // @[Cat.scala 29:58]
  wire [7:0] _GEN_172 = 10'hac == _T_7[9:0] ? 8'h13 : _GEN_171; // @[Cat.scala 29:58]
  wire [7:0] _GEN_173 = 10'had == _T_7[9:0] ? 8'h1 : _GEN_172; // @[Cat.scala 29:58]
  wire [7:0] _GEN_174 = 10'hae == _T_7[9:0] ? 8'h1 : _GEN_173; // @[Cat.scala 29:58]
  wire [7:0] _GEN_175 = 10'haf == _T_7[9:0] ? 8'hfe : _GEN_174; // @[Cat.scala 29:58]
  wire [7:0] _GEN_176 = 10'hb0 == _T_7[9:0] ? 8'h23 : _GEN_175; // @[Cat.scala 29:58]
  wire [7:0] _GEN_177 = 10'hb1 == _T_7[9:0] ? 8'h2e : _GEN_176; // @[Cat.scala 29:58]
  wire [7:0] _GEN_178 = 10'hb2 == _T_7[9:0] ? 8'h11 : _GEN_177; // @[Cat.scala 29:58]
  wire [7:0] _GEN_179 = 10'hb3 == _T_7[9:0] ? 8'h0 : _GEN_178; // @[Cat.scala 29:58]
  wire [7:0] _GEN_180 = 10'hb4 == _T_7[9:0] ? 8'h23 : _GEN_179; // @[Cat.scala 29:58]
  wire [7:0] _GEN_181 = 10'hb5 == _T_7[9:0] ? 8'h2c : _GEN_180; // @[Cat.scala 29:58]
  wire [7:0] _GEN_182 = 10'hb6 == _T_7[9:0] ? 8'h81 : _GEN_181; // @[Cat.scala 29:58]
  wire [7:0] _GEN_183 = 10'hb7 == _T_7[9:0] ? 8'h0 : _GEN_182; // @[Cat.scala 29:58]
  wire [7:0] _GEN_184 = 10'hb8 == _T_7[9:0] ? 8'h13 : _GEN_183; // @[Cat.scala 29:58]
  wire [7:0] _GEN_185 = 10'hb9 == _T_7[9:0] ? 8'h4 : _GEN_184; // @[Cat.scala 29:58]
  wire [7:0] _GEN_186 = 10'hba == _T_7[9:0] ? 8'h1 : _GEN_185; // @[Cat.scala 29:58]
  wire [7:0] _GEN_187 = 10'hbb == _T_7[9:0] ? 8'h2 : _GEN_186; // @[Cat.scala 29:58]
  wire [7:0] _GEN_188 = 10'hbc == _T_7[9:0] ? 8'h23 : _GEN_187; // @[Cat.scala 29:58]
  wire [7:0] _GEN_189 = 10'hbd == _T_7[9:0] ? 8'h26 : _GEN_188; // @[Cat.scala 29:58]
  wire [7:0] _GEN_190 = 10'hbe == _T_7[9:0] ? 8'h4 : _GEN_189; // @[Cat.scala 29:58]
  wire [7:0] _GEN_191 = 10'hbf == _T_7[9:0] ? 8'hfe : _GEN_190; // @[Cat.scala 29:58]
  wire [7:0] _GEN_192 = 10'hc0 == _T_7[9:0] ? 8'hb7 : _GEN_191; // @[Cat.scala 29:58]
  wire [7:0] _GEN_193 = 10'hc1 == _T_7[9:0] ? 8'hc7 : _GEN_192; // @[Cat.scala 29:58]
  wire [7:0] _GEN_194 = 10'hc2 == _T_7[9:0] ? 8'h0 : _GEN_193; // @[Cat.scala 29:58]
  wire [7:0] _GEN_195 = 10'hc3 == _T_7[9:0] ? 8'h0 : _GEN_194; // @[Cat.scala 29:58]
  wire [7:0] _GEN_196 = 10'hc4 == _T_7[9:0] ? 8'h13 : _GEN_195; // @[Cat.scala 29:58]
  wire [7:0] _GEN_197 = 10'hc5 == _T_7[9:0] ? 8'h85 : _GEN_196; // @[Cat.scala 29:58]
  wire [7:0] _GEN_198 = 10'hc6 == _T_7[9:0] ? 8'hf7 : _GEN_197; // @[Cat.scala 29:58]
  wire [7:0] _GEN_199 = 10'hc7 == _T_7[9:0] ? 8'hee : _GEN_198; // @[Cat.scala 29:58]
  wire [7:0] _GEN_200 = 10'hc8 == _T_7[9:0] ? 8'hef : _GEN_199; // @[Cat.scala 29:58]
  wire [7:0] _GEN_201 = 10'hc9 == _T_7[9:0] ? 8'hf0 : _GEN_200; // @[Cat.scala 29:58]
  wire [7:0] _GEN_202 = 10'hca == _T_7[9:0] ? 8'h1f : _GEN_201; // @[Cat.scala 29:58]
  wire [7:0] _GEN_203 = 10'hcb == _T_7[9:0] ? 8'hfb : _GEN_202; // @[Cat.scala 29:58]
  wire [7:0] _GEN_204 = 10'hcc == _T_7[9:0] ? 8'h23 : _GEN_203; // @[Cat.scala 29:58]
  wire [7:0] _GEN_205 = 10'hcd == _T_7[9:0] ? 8'h26 : _GEN_204; // @[Cat.scala 29:58]
  wire [7:0] _GEN_206 = 10'hce == _T_7[9:0] ? 8'h4 : _GEN_205; // @[Cat.scala 29:58]
  wire [7:0] _GEN_207 = 10'hcf == _T_7[9:0] ? 8'hfe : _GEN_206; // @[Cat.scala 29:58]
  wire [7:0] _GEN_208 = 10'hd0 == _T_7[9:0] ? 8'h6f : _GEN_207; // @[Cat.scala 29:58]
  wire [7:0] _GEN_209 = 10'hd1 == _T_7[9:0] ? 8'h0 : _GEN_208; // @[Cat.scala 29:58]
  wire [7:0] _GEN_210 = 10'hd2 == _T_7[9:0] ? 8'h0 : _GEN_209; // @[Cat.scala 29:58]
  wire [7:0] _GEN_211 = 10'hd3 == _T_7[9:0] ? 8'h1 : _GEN_210; // @[Cat.scala 29:58]
  wire [7:0] _GEN_212 = 10'hd4 == _T_7[9:0] ? 8'h83 : _GEN_211; // @[Cat.scala 29:58]
  wire [7:0] _GEN_213 = 10'hd5 == _T_7[9:0] ? 8'h27 : _GEN_212; // @[Cat.scala 29:58]
  wire [7:0] _GEN_214 = 10'hd6 == _T_7[9:0] ? 8'hc4 : _GEN_213; // @[Cat.scala 29:58]
  wire [7:0] _GEN_215 = 10'hd7 == _T_7[9:0] ? 8'hfe : _GEN_214; // @[Cat.scala 29:58]
  wire [7:0] _GEN_216 = 10'hd8 == _T_7[9:0] ? 8'h93 : _GEN_215; // @[Cat.scala 29:58]
  wire [7:0] _GEN_217 = 10'hd9 == _T_7[9:0] ? 8'h87 : _GEN_216; // @[Cat.scala 29:58]
  wire [7:0] _GEN_218 = 10'hda == _T_7[9:0] ? 8'h17 : _GEN_217; // @[Cat.scala 29:58]
  wire [7:0] _GEN_219 = 10'hdb == _T_7[9:0] ? 8'h0 : _GEN_218; // @[Cat.scala 29:58]
  wire [7:0] _GEN_220 = 10'hdc == _T_7[9:0] ? 8'h23 : _GEN_219; // @[Cat.scala 29:58]
  wire [7:0] _GEN_221 = 10'hdd == _T_7[9:0] ? 8'h26 : _GEN_220; // @[Cat.scala 29:58]
  wire [7:0] _GEN_222 = 10'hde == _T_7[9:0] ? 8'hf4 : _GEN_221; // @[Cat.scala 29:58]
  wire [7:0] _GEN_223 = 10'hdf == _T_7[9:0] ? 8'hfe : _GEN_222; // @[Cat.scala 29:58]
  wire [7:0] _GEN_224 = 10'he0 == _T_7[9:0] ? 8'h3 : _GEN_223; // @[Cat.scala 29:58]
  wire [7:0] _GEN_225 = 10'he1 == _T_7[9:0] ? 8'h27 : _GEN_224; // @[Cat.scala 29:58]
  wire [7:0] _GEN_226 = 10'he2 == _T_7[9:0] ? 8'hc4 : _GEN_225; // @[Cat.scala 29:58]
  wire [7:0] _GEN_227 = 10'he3 == _T_7[9:0] ? 8'hfe : _GEN_226; // @[Cat.scala 29:58]
  wire [7:0] _GEN_228 = 10'he4 == _T_7[9:0] ? 8'hb7 : _GEN_227; // @[Cat.scala 29:58]
  wire [7:0] _GEN_229 = 10'he5 == _T_7[9:0] ? 8'h17 : _GEN_228; // @[Cat.scala 29:58]
  wire [7:0] _GEN_230 = 10'he6 == _T_7[9:0] ? 8'h7a : _GEN_229; // @[Cat.scala 29:58]
  wire [7:0] _GEN_231 = 10'he7 == _T_7[9:0] ? 8'h0 : _GEN_230; // @[Cat.scala 29:58]
  wire [7:0] _GEN_232 = 10'he8 == _T_7[9:0] ? 8'h93 : _GEN_231; // @[Cat.scala 29:58]
  wire [7:0] _GEN_233 = 10'he9 == _T_7[9:0] ? 8'h87 : _GEN_232; // @[Cat.scala 29:58]
  wire [7:0] _GEN_234 = 10'hea == _T_7[9:0] ? 8'hf7 : _GEN_233; // @[Cat.scala 29:58]
  wire [7:0] _GEN_235 = 10'heb == _T_7[9:0] ? 8'h1f : _GEN_234; // @[Cat.scala 29:58]
  wire [7:0] _GEN_236 = 10'hec == _T_7[9:0] ? 8'he3 : _GEN_235; // @[Cat.scala 29:58]
  wire [7:0] _GEN_237 = 10'hed == _T_7[9:0] ? 8'hd4 : _GEN_236; // @[Cat.scala 29:58]
  wire [7:0] _GEN_238 = 10'hee == _T_7[9:0] ? 8'he7 : _GEN_237; // @[Cat.scala 29:58]
  wire [7:0] _GEN_239 = 10'hef == _T_7[9:0] ? 8'hfe : _GEN_238; // @[Cat.scala 29:58]
  wire [7:0] _GEN_240 = 10'hf0 == _T_7[9:0] ? 8'h13 : _GEN_239; // @[Cat.scala 29:58]
  wire [7:0] _GEN_241 = 10'hf1 == _T_7[9:0] ? 8'h5 : _GEN_240; // @[Cat.scala 29:58]
  wire [7:0] _GEN_242 = 10'hf2 == _T_7[9:0] ? 8'h0 : _GEN_241; // @[Cat.scala 29:58]
  wire [7:0] _GEN_243 = 10'hf3 == _T_7[9:0] ? 8'h0 : _GEN_242; // @[Cat.scala 29:58]
  wire [7:0] _GEN_244 = 10'hf4 == _T_7[9:0] ? 8'hef : _GEN_243; // @[Cat.scala 29:58]
  wire [7:0] _GEN_245 = 10'hf5 == _T_7[9:0] ? 8'hf0 : _GEN_244; // @[Cat.scala 29:58]
  wire [7:0] _GEN_246 = 10'hf6 == _T_7[9:0] ? 8'h5f : _GEN_245; // @[Cat.scala 29:58]
  wire [7:0] _GEN_247 = 10'hf7 == _T_7[9:0] ? 8'hf8 : _GEN_246; // @[Cat.scala 29:58]
  wire [7:0] _GEN_248 = 10'hf8 == _T_7[9:0] ? 8'hef : _GEN_247; // @[Cat.scala 29:58]
  wire [7:0] _GEN_249 = 10'hf9 == _T_7[9:0] ? 8'hf0 : _GEN_248; // @[Cat.scala 29:58]
  wire [7:0] _GEN_250 = 10'hfa == _T_7[9:0] ? 8'h1f : _GEN_249; // @[Cat.scala 29:58]
  wire [7:0] _GEN_251 = 10'hfb == _T_7[9:0] ? 8'hf5 : _GEN_250; // @[Cat.scala 29:58]
  wire [7:0] _GEN_252 = 10'hfc == _T_7[9:0] ? 8'h93 : _GEN_251; // @[Cat.scala 29:58]
  wire [7:0] _GEN_253 = 10'hfd == _T_7[9:0] ? 8'h7 : _GEN_252; // @[Cat.scala 29:58]
  wire [7:0] _GEN_254 = 10'hfe == _T_7[9:0] ? 8'h5 : _GEN_253; // @[Cat.scala 29:58]
  wire [7:0] _GEN_255 = 10'hff == _T_7[9:0] ? 8'h0 : _GEN_254; // @[Cat.scala 29:58]
  wire [7:0] _GEN_256 = 10'h100 == _T_7[9:0] ? 8'he3 : _GEN_255; // @[Cat.scala 29:58]
  wire [7:0] _GEN_257 = 10'h101 == _T_7[9:0] ? 8'h8c : _GEN_256; // @[Cat.scala 29:58]
  wire [7:0] _GEN_258 = 10'h102 == _T_7[9:0] ? 8'h7 : _GEN_257; // @[Cat.scala 29:58]
  wire [7:0] _GEN_259 = 10'h103 == _T_7[9:0] ? 8'hfe : _GEN_258; // @[Cat.scala 29:58]
  wire [7:0] _GEN_260 = 10'h104 == _T_7[9:0] ? 8'hef : _GEN_259; // @[Cat.scala 29:58]
  wire [7:0] _GEN_261 = 10'h105 == _T_7[9:0] ? 8'hf0 : _GEN_260; // @[Cat.scala 29:58]
  wire [7:0] _GEN_262 = 10'h106 == _T_7[9:0] ? 8'h5f : _GEN_261; // @[Cat.scala 29:58]
  wire [7:0] _GEN_263 = 10'h107 == _T_7[9:0] ? 8'hf1 : _GEN_262; // @[Cat.scala 29:58]
  wire [7:0] _GEN_264 = 10'h108 == _T_7[9:0] ? 8'h93 : _GEN_263; // @[Cat.scala 29:58]
  wire [7:0] _GEN_265 = 10'h109 == _T_7[9:0] ? 8'h7 : _GEN_264; // @[Cat.scala 29:58]
  wire [7:0] _GEN_266 = 10'h10a == _T_7[9:0] ? 8'h5 : _GEN_265; // @[Cat.scala 29:58]
  wire [7:0] _GEN_267 = 10'h10b == _T_7[9:0] ? 8'h0 : _GEN_266; // @[Cat.scala 29:58]
  wire [7:0] _GEN_268 = 10'h10c == _T_7[9:0] ? 8'h13 : _GEN_267; // @[Cat.scala 29:58]
  wire [7:0] _GEN_269 = 10'h10d == _T_7[9:0] ? 8'h85 : _GEN_268; // @[Cat.scala 29:58]
  wire [7:0] _GEN_270 = 10'h10e == _T_7[9:0] ? 8'h7 : _GEN_269; // @[Cat.scala 29:58]
  wire [7:0] _GEN_271 = 10'h10f == _T_7[9:0] ? 8'h0 : _GEN_270; // @[Cat.scala 29:58]
  wire [7:0] _GEN_272 = 10'h110 == _T_7[9:0] ? 8'hef : _GEN_271; // @[Cat.scala 29:58]
  wire [7:0] _GEN_273 = 10'h111 == _T_7[9:0] ? 8'hf0 : _GEN_272; // @[Cat.scala 29:58]
  wire [7:0] _GEN_274 = 10'h112 == _T_7[9:0] ? 8'h9f : _GEN_273; // @[Cat.scala 29:58]
  wire [7:0] _GEN_275 = 10'h113 == _T_7[9:0] ? 8'hf6 : _GEN_274; // @[Cat.scala 29:58]
  wire [7:0] _GEN_276 = 10'h114 == _T_7[9:0] ? 8'h23 : _GEN_275; // @[Cat.scala 29:58]
  wire [7:0] _GEN_277 = 10'h115 == _T_7[9:0] ? 8'h26 : _GEN_276; // @[Cat.scala 29:58]
  wire [7:0] _GEN_278 = 10'h116 == _T_7[9:0] ? 8'h4 : _GEN_277; // @[Cat.scala 29:58]
  wire [7:0] _GEN_279 = 10'h117 == _T_7[9:0] ? 8'hfe : _GEN_278; // @[Cat.scala 29:58]
  wire [7:0] _GEN_280 = 10'h118 == _T_7[9:0] ? 8'h6f : _GEN_279; // @[Cat.scala 29:58]
  wire [7:0] _GEN_281 = 10'h119 == _T_7[9:0] ? 8'h0 : _GEN_280; // @[Cat.scala 29:58]
  wire [7:0] _GEN_282 = 10'h11a == _T_7[9:0] ? 8'h0 : _GEN_281; // @[Cat.scala 29:58]
  wire [7:0] _GEN_283 = 10'h11b == _T_7[9:0] ? 8'h1 : _GEN_282; // @[Cat.scala 29:58]
  wire [7:0] _GEN_284 = 10'h11c == _T_7[9:0] ? 8'h83 : _GEN_283; // @[Cat.scala 29:58]
  wire [7:0] _GEN_285 = 10'h11d == _T_7[9:0] ? 8'h27 : _GEN_284; // @[Cat.scala 29:58]
  wire [7:0] _GEN_286 = 10'h11e == _T_7[9:0] ? 8'hc4 : _GEN_285; // @[Cat.scala 29:58]
  wire [7:0] _GEN_287 = 10'h11f == _T_7[9:0] ? 8'hfe : _GEN_286; // @[Cat.scala 29:58]
  wire [7:0] _GEN_288 = 10'h120 == _T_7[9:0] ? 8'h93 : _GEN_287; // @[Cat.scala 29:58]
  wire [7:0] _GEN_289 = 10'h121 == _T_7[9:0] ? 8'h87 : _GEN_288; // @[Cat.scala 29:58]
  wire [7:0] _GEN_290 = 10'h122 == _T_7[9:0] ? 8'h17 : _GEN_289; // @[Cat.scala 29:58]
  wire [7:0] _GEN_291 = 10'h123 == _T_7[9:0] ? 8'h0 : _GEN_290; // @[Cat.scala 29:58]
  wire [7:0] _GEN_292 = 10'h124 == _T_7[9:0] ? 8'h23 : _GEN_291; // @[Cat.scala 29:58]
  wire [7:0] _GEN_293 = 10'h125 == _T_7[9:0] ? 8'h26 : _GEN_292; // @[Cat.scala 29:58]
  wire [7:0] _GEN_294 = 10'h126 == _T_7[9:0] ? 8'hf4 : _GEN_293; // @[Cat.scala 29:58]
  wire [7:0] _GEN_295 = 10'h127 == _T_7[9:0] ? 8'hfe : _GEN_294; // @[Cat.scala 29:58]
  wire [7:0] _GEN_296 = 10'h128 == _T_7[9:0] ? 8'h3 : _GEN_295; // @[Cat.scala 29:58]
  wire [7:0] _GEN_297 = 10'h129 == _T_7[9:0] ? 8'h27 : _GEN_296; // @[Cat.scala 29:58]
  wire [7:0] _GEN_298 = 10'h12a == _T_7[9:0] ? 8'hc4 : _GEN_297; // @[Cat.scala 29:58]
  wire [7:0] _GEN_299 = 10'h12b == _T_7[9:0] ? 8'hfe : _GEN_298; // @[Cat.scala 29:58]
  wire [7:0] _GEN_300 = 10'h12c == _T_7[9:0] ? 8'hb7 : _GEN_299; // @[Cat.scala 29:58]
  wire [7:0] _GEN_301 = 10'h12d == _T_7[9:0] ? 8'h57 : _GEN_300; // @[Cat.scala 29:58]
  wire [7:0] _GEN_302 = 10'h12e == _T_7[9:0] ? 8'h89 : _GEN_301; // @[Cat.scala 29:58]
  wire [7:0] _GEN_303 = 10'h12f == _T_7[9:0] ? 8'h0 : _GEN_302; // @[Cat.scala 29:58]
  wire [7:0] _GEN_304 = 10'h130 == _T_7[9:0] ? 8'h93 : _GEN_303; // @[Cat.scala 29:58]
  wire [7:0] _GEN_305 = 10'h131 == _T_7[9:0] ? 8'h87 : _GEN_304; // @[Cat.scala 29:58]
  wire [7:0] _GEN_306 = 10'h132 == _T_7[9:0] ? 8'hf7 : _GEN_305; // @[Cat.scala 29:58]
  wire [7:0] _GEN_307 = 10'h133 == _T_7[9:0] ? 8'h43 : _GEN_306; // @[Cat.scala 29:58]
  wire [7:0] _GEN_308 = 10'h134 == _T_7[9:0] ? 8'he3 : _GEN_307; // @[Cat.scala 29:58]
  wire [7:0] _GEN_309 = 10'h135 == _T_7[9:0] ? 8'hd4 : _GEN_308; // @[Cat.scala 29:58]
  wire [7:0] _GEN_310 = 10'h136 == _T_7[9:0] ? 8'he7 : _GEN_309; // @[Cat.scala 29:58]
  wire [7:0] _GEN_311 = 10'h137 == _T_7[9:0] ? 8'hfe : _GEN_310; // @[Cat.scala 29:58]
  wire [7:0] _GEN_312 = 10'h138 == _T_7[9:0] ? 8'h13 : _GEN_311; // @[Cat.scala 29:58]
  wire [7:0] _GEN_313 = 10'h139 == _T_7[9:0] ? 8'h5 : _GEN_312; // @[Cat.scala 29:58]
  wire [7:0] _GEN_314 = 10'h13a == _T_7[9:0] ? 8'h0 : _GEN_313; // @[Cat.scala 29:58]
  wire [7:0] _GEN_315 = 10'h13b == _T_7[9:0] ? 8'h0 : _GEN_314; // @[Cat.scala 29:58]
  wire [7:0] _GEN_316 = 10'h13c == _T_7[9:0] ? 8'hef : _GEN_315; // @[Cat.scala 29:58]
  wire [7:0] _GEN_317 = 10'h13d == _T_7[9:0] ? 8'hf0 : _GEN_316; // @[Cat.scala 29:58]
  wire [7:0] _GEN_318 = 10'h13e == _T_7[9:0] ? 8'hdf : _GEN_317; // @[Cat.scala 29:58]
  wire [7:0] _GEN_319 = 10'h13f == _T_7[9:0] ? 8'hf3 : _GEN_318; // @[Cat.scala 29:58]
  wire [7:0] _GEN_320 = 10'h140 == _T_7[9:0] ? 8'h6f : _GEN_319; // @[Cat.scala 29:58]
  wire [7:0] _GEN_321 = 10'h141 == _T_7[9:0] ? 8'hf0 : _GEN_320; // @[Cat.scala 29:58]
  wire [7:0] _GEN_322 = 10'h142 == _T_7[9:0] ? 8'h9f : _GEN_321; // @[Cat.scala 29:58]
  wire [7:0] _GEN_323 = 10'h143 == _T_7[9:0] ? 8'hfb : _GEN_322; // @[Cat.scala 29:58]
  wire [7:0] _GEN_324 = 10'h144 == _T_7[9:0] ? 8'h0 : _GEN_323; // @[Cat.scala 29:58]
  wire [7:0] _GEN_325 = 10'h145 == _T_7[9:0] ? 8'h0 : _GEN_324; // @[Cat.scala 29:58]
  wire [7:0] _GEN_326 = 10'h146 == _T_7[9:0] ? 8'h0 : _GEN_325; // @[Cat.scala 29:58]
  wire [7:0] _GEN_327 = 10'h147 == _T_7[9:0] ? 8'h0 : _GEN_326; // @[Cat.scala 29:58]
  wire [7:0] _GEN_328 = 10'h148 == _T_7[9:0] ? 8'h0 : _GEN_327; // @[Cat.scala 29:58]
  wire [7:0] _GEN_329 = 10'h149 == _T_7[9:0] ? 8'h0 : _GEN_328; // @[Cat.scala 29:58]
  wire [7:0] _GEN_330 = 10'h14a == _T_7[9:0] ? 8'h0 : _GEN_329; // @[Cat.scala 29:58]
  wire [7:0] _GEN_331 = 10'h14b == _T_7[9:0] ? 8'h0 : _GEN_330; // @[Cat.scala 29:58]
  wire [7:0] _GEN_332 = 10'h14c == _T_7[9:0] ? 8'h0 : _GEN_331; // @[Cat.scala 29:58]
  wire [7:0] _GEN_333 = 10'h14d == _T_7[9:0] ? 8'h0 : _GEN_332; // @[Cat.scala 29:58]
  wire [7:0] _GEN_334 = 10'h14e == _T_7[9:0] ? 8'h0 : _GEN_333; // @[Cat.scala 29:58]
  wire [7:0] _GEN_335 = 10'h14f == _T_7[9:0] ? 8'h0 : _GEN_334; // @[Cat.scala 29:58]
  wire [7:0] _GEN_336 = 10'h150 == _T_7[9:0] ? 8'h0 : _GEN_335; // @[Cat.scala 29:58]
  wire [7:0] _GEN_337 = 10'h151 == _T_7[9:0] ? 8'h0 : _GEN_336; // @[Cat.scala 29:58]
  wire [7:0] _GEN_338 = 10'h152 == _T_7[9:0] ? 8'h0 : _GEN_337; // @[Cat.scala 29:58]
  wire [7:0] _GEN_339 = 10'h153 == _T_7[9:0] ? 8'h0 : _GEN_338; // @[Cat.scala 29:58]
  wire [7:0] _GEN_340 = 10'h154 == _T_7[9:0] ? 8'h0 : _GEN_339; // @[Cat.scala 29:58]
  wire [7:0] _GEN_341 = 10'h155 == _T_7[9:0] ? 8'h0 : _GEN_340; // @[Cat.scala 29:58]
  wire [7:0] _GEN_342 = 10'h156 == _T_7[9:0] ? 8'h0 : _GEN_341; // @[Cat.scala 29:58]
  wire [7:0] _GEN_343 = 10'h157 == _T_7[9:0] ? 8'h0 : _GEN_342; // @[Cat.scala 29:58]
  wire [7:0] _GEN_344 = 10'h158 == _T_7[9:0] ? 8'h0 : _GEN_343; // @[Cat.scala 29:58]
  wire [7:0] _GEN_345 = 10'h159 == _T_7[9:0] ? 8'h0 : _GEN_344; // @[Cat.scala 29:58]
  wire [7:0] _GEN_346 = 10'h15a == _T_7[9:0] ? 8'h0 : _GEN_345; // @[Cat.scala 29:58]
  wire [7:0] _GEN_347 = 10'h15b == _T_7[9:0] ? 8'h0 : _GEN_346; // @[Cat.scala 29:58]
  wire [7:0] _GEN_348 = 10'h15c == _T_7[9:0] ? 8'h0 : _GEN_347; // @[Cat.scala 29:58]
  wire [7:0] _GEN_349 = 10'h15d == _T_7[9:0] ? 8'h0 : _GEN_348; // @[Cat.scala 29:58]
  wire [7:0] _GEN_350 = 10'h15e == _T_7[9:0] ? 8'h0 : _GEN_349; // @[Cat.scala 29:58]
  wire [7:0] _GEN_351 = 10'h15f == _T_7[9:0] ? 8'h0 : _GEN_350; // @[Cat.scala 29:58]
  wire [7:0] _GEN_352 = 10'h160 == _T_7[9:0] ? 8'h0 : _GEN_351; // @[Cat.scala 29:58]
  wire [7:0] _GEN_353 = 10'h161 == _T_7[9:0] ? 8'h0 : _GEN_352; // @[Cat.scala 29:58]
  wire [7:0] _GEN_354 = 10'h162 == _T_7[9:0] ? 8'h0 : _GEN_353; // @[Cat.scala 29:58]
  wire [7:0] _GEN_355 = 10'h163 == _T_7[9:0] ? 8'h0 : _GEN_354; // @[Cat.scala 29:58]
  wire [7:0] _GEN_356 = 10'h164 == _T_7[9:0] ? 8'h0 : _GEN_355; // @[Cat.scala 29:58]
  wire [7:0] _GEN_357 = 10'h165 == _T_7[9:0] ? 8'h0 : _GEN_356; // @[Cat.scala 29:58]
  wire [7:0] _GEN_358 = 10'h166 == _T_7[9:0] ? 8'h0 : _GEN_357; // @[Cat.scala 29:58]
  wire [7:0] _GEN_359 = 10'h167 == _T_7[9:0] ? 8'h0 : _GEN_358; // @[Cat.scala 29:58]
  wire [7:0] _GEN_360 = 10'h168 == _T_7[9:0] ? 8'h0 : _GEN_359; // @[Cat.scala 29:58]
  wire [7:0] _GEN_361 = 10'h169 == _T_7[9:0] ? 8'h0 : _GEN_360; // @[Cat.scala 29:58]
  wire [7:0] _GEN_362 = 10'h16a == _T_7[9:0] ? 8'h0 : _GEN_361; // @[Cat.scala 29:58]
  wire [7:0] _GEN_363 = 10'h16b == _T_7[9:0] ? 8'h0 : _GEN_362; // @[Cat.scala 29:58]
  wire [7:0] _GEN_364 = 10'h16c == _T_7[9:0] ? 8'h0 : _GEN_363; // @[Cat.scala 29:58]
  wire [7:0] _GEN_365 = 10'h16d == _T_7[9:0] ? 8'h0 : _GEN_364; // @[Cat.scala 29:58]
  wire [7:0] _GEN_366 = 10'h16e == _T_7[9:0] ? 8'h0 : _GEN_365; // @[Cat.scala 29:58]
  wire [7:0] _GEN_367 = 10'h16f == _T_7[9:0] ? 8'h0 : _GEN_366; // @[Cat.scala 29:58]
  wire [7:0] _GEN_368 = 10'h170 == _T_7[9:0] ? 8'h0 : _GEN_367; // @[Cat.scala 29:58]
  wire [7:0] _GEN_369 = 10'h171 == _T_7[9:0] ? 8'h0 : _GEN_368; // @[Cat.scala 29:58]
  wire [7:0] _GEN_370 = 10'h172 == _T_7[9:0] ? 8'h0 : _GEN_369; // @[Cat.scala 29:58]
  wire [7:0] _GEN_371 = 10'h173 == _T_7[9:0] ? 8'h0 : _GEN_370; // @[Cat.scala 29:58]
  wire [7:0] _GEN_372 = 10'h174 == _T_7[9:0] ? 8'h0 : _GEN_371; // @[Cat.scala 29:58]
  wire [7:0] _GEN_373 = 10'h175 == _T_7[9:0] ? 8'h0 : _GEN_372; // @[Cat.scala 29:58]
  wire [7:0] _GEN_374 = 10'h176 == _T_7[9:0] ? 8'h0 : _GEN_373; // @[Cat.scala 29:58]
  wire [7:0] _GEN_375 = 10'h177 == _T_7[9:0] ? 8'h0 : _GEN_374; // @[Cat.scala 29:58]
  wire [7:0] _GEN_376 = 10'h178 == _T_7[9:0] ? 8'h0 : _GEN_375; // @[Cat.scala 29:58]
  wire [7:0] _GEN_377 = 10'h179 == _T_7[9:0] ? 8'h0 : _GEN_376; // @[Cat.scala 29:58]
  wire [7:0] _GEN_378 = 10'h17a == _T_7[9:0] ? 8'h0 : _GEN_377; // @[Cat.scala 29:58]
  wire [7:0] _GEN_379 = 10'h17b == _T_7[9:0] ? 8'h0 : _GEN_378; // @[Cat.scala 29:58]
  wire [7:0] _GEN_380 = 10'h17c == _T_7[9:0] ? 8'h0 : _GEN_379; // @[Cat.scala 29:58]
  wire [7:0] _GEN_381 = 10'h17d == _T_7[9:0] ? 8'h0 : _GEN_380; // @[Cat.scala 29:58]
  wire [7:0] _GEN_382 = 10'h17e == _T_7[9:0] ? 8'h0 : _GEN_381; // @[Cat.scala 29:58]
  wire [7:0] _GEN_383 = 10'h17f == _T_7[9:0] ? 8'h0 : _GEN_382; // @[Cat.scala 29:58]
  wire [7:0] _GEN_384 = 10'h180 == _T_7[9:0] ? 8'h0 : _GEN_383; // @[Cat.scala 29:58]
  wire [7:0] _GEN_385 = 10'h181 == _T_7[9:0] ? 8'h0 : _GEN_384; // @[Cat.scala 29:58]
  wire [7:0] _GEN_386 = 10'h182 == _T_7[9:0] ? 8'h0 : _GEN_385; // @[Cat.scala 29:58]
  wire [7:0] _GEN_387 = 10'h183 == _T_7[9:0] ? 8'h0 : _GEN_386; // @[Cat.scala 29:58]
  wire [7:0] _GEN_388 = 10'h184 == _T_7[9:0] ? 8'h0 : _GEN_387; // @[Cat.scala 29:58]
  wire [7:0] _GEN_389 = 10'h185 == _T_7[9:0] ? 8'h0 : _GEN_388; // @[Cat.scala 29:58]
  wire [7:0] _GEN_390 = 10'h186 == _T_7[9:0] ? 8'h0 : _GEN_389; // @[Cat.scala 29:58]
  wire [7:0] _GEN_391 = 10'h187 == _T_7[9:0] ? 8'h0 : _GEN_390; // @[Cat.scala 29:58]
  wire [7:0] _GEN_392 = 10'h188 == _T_7[9:0] ? 8'h0 : _GEN_391; // @[Cat.scala 29:58]
  wire [7:0] _GEN_393 = 10'h189 == _T_7[9:0] ? 8'h0 : _GEN_392; // @[Cat.scala 29:58]
  wire [7:0] _GEN_394 = 10'h18a == _T_7[9:0] ? 8'h0 : _GEN_393; // @[Cat.scala 29:58]
  wire [7:0] _GEN_395 = 10'h18b == _T_7[9:0] ? 8'h0 : _GEN_394; // @[Cat.scala 29:58]
  wire [7:0] _GEN_396 = 10'h18c == _T_7[9:0] ? 8'h0 : _GEN_395; // @[Cat.scala 29:58]
  wire [7:0] _GEN_397 = 10'h18d == _T_7[9:0] ? 8'h0 : _GEN_396; // @[Cat.scala 29:58]
  wire [7:0] _GEN_398 = 10'h18e == _T_7[9:0] ? 8'h0 : _GEN_397; // @[Cat.scala 29:58]
  wire [7:0] _GEN_399 = 10'h18f == _T_7[9:0] ? 8'h0 : _GEN_398; // @[Cat.scala 29:58]
  wire [7:0] _GEN_400 = 10'h190 == _T_7[9:0] ? 8'h0 : _GEN_399; // @[Cat.scala 29:58]
  wire [7:0] _GEN_401 = 10'h191 == _T_7[9:0] ? 8'h0 : _GEN_400; // @[Cat.scala 29:58]
  wire [7:0] _GEN_402 = 10'h192 == _T_7[9:0] ? 8'h0 : _GEN_401; // @[Cat.scala 29:58]
  wire [7:0] _GEN_403 = 10'h193 == _T_7[9:0] ? 8'h0 : _GEN_402; // @[Cat.scala 29:58]
  wire [7:0] _GEN_404 = 10'h194 == _T_7[9:0] ? 8'h0 : _GEN_403; // @[Cat.scala 29:58]
  wire [7:0] _GEN_405 = 10'h195 == _T_7[9:0] ? 8'h0 : _GEN_404; // @[Cat.scala 29:58]
  wire [7:0] _GEN_406 = 10'h196 == _T_7[9:0] ? 8'h0 : _GEN_405; // @[Cat.scala 29:58]
  wire [7:0] _GEN_407 = 10'h197 == _T_7[9:0] ? 8'h0 : _GEN_406; // @[Cat.scala 29:58]
  wire [7:0] _GEN_408 = 10'h198 == _T_7[9:0] ? 8'h0 : _GEN_407; // @[Cat.scala 29:58]
  wire [7:0] _GEN_409 = 10'h199 == _T_7[9:0] ? 8'h0 : _GEN_408; // @[Cat.scala 29:58]
  wire [7:0] _GEN_410 = 10'h19a == _T_7[9:0] ? 8'h0 : _GEN_409; // @[Cat.scala 29:58]
  wire [7:0] _GEN_411 = 10'h19b == _T_7[9:0] ? 8'h0 : _GEN_410; // @[Cat.scala 29:58]
  wire [7:0] _GEN_412 = 10'h19c == _T_7[9:0] ? 8'h0 : _GEN_411; // @[Cat.scala 29:58]
  wire [7:0] _GEN_413 = 10'h19d == _T_7[9:0] ? 8'h0 : _GEN_412; // @[Cat.scala 29:58]
  wire [7:0] _GEN_414 = 10'h19e == _T_7[9:0] ? 8'h0 : _GEN_413; // @[Cat.scala 29:58]
  wire [7:0] _GEN_415 = 10'h19f == _T_7[9:0] ? 8'h0 : _GEN_414; // @[Cat.scala 29:58]
  wire [7:0] _GEN_416 = 10'h1a0 == _T_7[9:0] ? 8'h0 : _GEN_415; // @[Cat.scala 29:58]
  wire [7:0] _GEN_417 = 10'h1a1 == _T_7[9:0] ? 8'h0 : _GEN_416; // @[Cat.scala 29:58]
  wire [7:0] _GEN_418 = 10'h1a2 == _T_7[9:0] ? 8'h0 : _GEN_417; // @[Cat.scala 29:58]
  wire [7:0] _GEN_419 = 10'h1a3 == _T_7[9:0] ? 8'h0 : _GEN_418; // @[Cat.scala 29:58]
  wire [7:0] _GEN_420 = 10'h1a4 == _T_7[9:0] ? 8'h0 : _GEN_419; // @[Cat.scala 29:58]
  wire [7:0] _GEN_421 = 10'h1a5 == _T_7[9:0] ? 8'h0 : _GEN_420; // @[Cat.scala 29:58]
  wire [7:0] _GEN_422 = 10'h1a6 == _T_7[9:0] ? 8'h0 : _GEN_421; // @[Cat.scala 29:58]
  wire [7:0] _GEN_423 = 10'h1a7 == _T_7[9:0] ? 8'h0 : _GEN_422; // @[Cat.scala 29:58]
  wire [7:0] _GEN_424 = 10'h1a8 == _T_7[9:0] ? 8'h0 : _GEN_423; // @[Cat.scala 29:58]
  wire [7:0] _GEN_425 = 10'h1a9 == _T_7[9:0] ? 8'h0 : _GEN_424; // @[Cat.scala 29:58]
  wire [7:0] _GEN_426 = 10'h1aa == _T_7[9:0] ? 8'h0 : _GEN_425; // @[Cat.scala 29:58]
  wire [7:0] _GEN_427 = 10'h1ab == _T_7[9:0] ? 8'h0 : _GEN_426; // @[Cat.scala 29:58]
  wire [7:0] _GEN_428 = 10'h1ac == _T_7[9:0] ? 8'h0 : _GEN_427; // @[Cat.scala 29:58]
  wire [7:0] _GEN_429 = 10'h1ad == _T_7[9:0] ? 8'h0 : _GEN_428; // @[Cat.scala 29:58]
  wire [7:0] _GEN_430 = 10'h1ae == _T_7[9:0] ? 8'h0 : _GEN_429; // @[Cat.scala 29:58]
  wire [7:0] _GEN_431 = 10'h1af == _T_7[9:0] ? 8'h0 : _GEN_430; // @[Cat.scala 29:58]
  wire [7:0] _GEN_432 = 10'h1b0 == _T_7[9:0] ? 8'h0 : _GEN_431; // @[Cat.scala 29:58]
  wire [7:0] _GEN_433 = 10'h1b1 == _T_7[9:0] ? 8'h0 : _GEN_432; // @[Cat.scala 29:58]
  wire [7:0] _GEN_434 = 10'h1b2 == _T_7[9:0] ? 8'h0 : _GEN_433; // @[Cat.scala 29:58]
  wire [7:0] _GEN_435 = 10'h1b3 == _T_7[9:0] ? 8'h0 : _GEN_434; // @[Cat.scala 29:58]
  wire [7:0] _GEN_436 = 10'h1b4 == _T_7[9:0] ? 8'h0 : _GEN_435; // @[Cat.scala 29:58]
  wire [7:0] _GEN_437 = 10'h1b5 == _T_7[9:0] ? 8'h0 : _GEN_436; // @[Cat.scala 29:58]
  wire [7:0] _GEN_438 = 10'h1b6 == _T_7[9:0] ? 8'h0 : _GEN_437; // @[Cat.scala 29:58]
  wire [7:0] _GEN_439 = 10'h1b7 == _T_7[9:0] ? 8'h0 : _GEN_438; // @[Cat.scala 29:58]
  wire [7:0] _GEN_440 = 10'h1b8 == _T_7[9:0] ? 8'h0 : _GEN_439; // @[Cat.scala 29:58]
  wire [7:0] _GEN_441 = 10'h1b9 == _T_7[9:0] ? 8'h0 : _GEN_440; // @[Cat.scala 29:58]
  wire [7:0] _GEN_442 = 10'h1ba == _T_7[9:0] ? 8'h0 : _GEN_441; // @[Cat.scala 29:58]
  wire [7:0] _GEN_443 = 10'h1bb == _T_7[9:0] ? 8'h0 : _GEN_442; // @[Cat.scala 29:58]
  wire [7:0] _GEN_444 = 10'h1bc == _T_7[9:0] ? 8'h0 : _GEN_443; // @[Cat.scala 29:58]
  wire [7:0] _GEN_445 = 10'h1bd == _T_7[9:0] ? 8'h0 : _GEN_444; // @[Cat.scala 29:58]
  wire [7:0] _GEN_446 = 10'h1be == _T_7[9:0] ? 8'h0 : _GEN_445; // @[Cat.scala 29:58]
  wire [7:0] _GEN_447 = 10'h1bf == _T_7[9:0] ? 8'h0 : _GEN_446; // @[Cat.scala 29:58]
  wire [7:0] _GEN_448 = 10'h1c0 == _T_7[9:0] ? 8'h0 : _GEN_447; // @[Cat.scala 29:58]
  wire [7:0] _GEN_449 = 10'h1c1 == _T_7[9:0] ? 8'h0 : _GEN_448; // @[Cat.scala 29:58]
  wire [7:0] _GEN_450 = 10'h1c2 == _T_7[9:0] ? 8'h0 : _GEN_449; // @[Cat.scala 29:58]
  wire [7:0] _GEN_451 = 10'h1c3 == _T_7[9:0] ? 8'h0 : _GEN_450; // @[Cat.scala 29:58]
  wire [7:0] _GEN_452 = 10'h1c4 == _T_7[9:0] ? 8'h0 : _GEN_451; // @[Cat.scala 29:58]
  wire [7:0] _GEN_453 = 10'h1c5 == _T_7[9:0] ? 8'h0 : _GEN_452; // @[Cat.scala 29:58]
  wire [7:0] _GEN_454 = 10'h1c6 == _T_7[9:0] ? 8'h0 : _GEN_453; // @[Cat.scala 29:58]
  wire [7:0] _GEN_455 = 10'h1c7 == _T_7[9:0] ? 8'h0 : _GEN_454; // @[Cat.scala 29:58]
  wire [7:0] _GEN_456 = 10'h1c8 == _T_7[9:0] ? 8'h0 : _GEN_455; // @[Cat.scala 29:58]
  wire [7:0] _GEN_457 = 10'h1c9 == _T_7[9:0] ? 8'h0 : _GEN_456; // @[Cat.scala 29:58]
  wire [7:0] _GEN_458 = 10'h1ca == _T_7[9:0] ? 8'h0 : _GEN_457; // @[Cat.scala 29:58]
  wire [7:0] _GEN_459 = 10'h1cb == _T_7[9:0] ? 8'h0 : _GEN_458; // @[Cat.scala 29:58]
  wire [7:0] _GEN_460 = 10'h1cc == _T_7[9:0] ? 8'h0 : _GEN_459; // @[Cat.scala 29:58]
  wire [7:0] _GEN_461 = 10'h1cd == _T_7[9:0] ? 8'h0 : _GEN_460; // @[Cat.scala 29:58]
  wire [7:0] _GEN_462 = 10'h1ce == _T_7[9:0] ? 8'h0 : _GEN_461; // @[Cat.scala 29:58]
  wire [7:0] _GEN_463 = 10'h1cf == _T_7[9:0] ? 8'h0 : _GEN_462; // @[Cat.scala 29:58]
  wire [7:0] _GEN_464 = 10'h1d0 == _T_7[9:0] ? 8'h0 : _GEN_463; // @[Cat.scala 29:58]
  wire [7:0] _GEN_465 = 10'h1d1 == _T_7[9:0] ? 8'h0 : _GEN_464; // @[Cat.scala 29:58]
  wire [7:0] _GEN_466 = 10'h1d2 == _T_7[9:0] ? 8'h0 : _GEN_465; // @[Cat.scala 29:58]
  wire [7:0] _GEN_467 = 10'h1d3 == _T_7[9:0] ? 8'h0 : _GEN_466; // @[Cat.scala 29:58]
  wire [7:0] _GEN_468 = 10'h1d4 == _T_7[9:0] ? 8'h0 : _GEN_467; // @[Cat.scala 29:58]
  wire [7:0] _GEN_469 = 10'h1d5 == _T_7[9:0] ? 8'h0 : _GEN_468; // @[Cat.scala 29:58]
  wire [7:0] _GEN_470 = 10'h1d6 == _T_7[9:0] ? 8'h0 : _GEN_469; // @[Cat.scala 29:58]
  wire [7:0] _GEN_471 = 10'h1d7 == _T_7[9:0] ? 8'h0 : _GEN_470; // @[Cat.scala 29:58]
  wire [7:0] _GEN_472 = 10'h1d8 == _T_7[9:0] ? 8'h0 : _GEN_471; // @[Cat.scala 29:58]
  wire [7:0] _GEN_473 = 10'h1d9 == _T_7[9:0] ? 8'h0 : _GEN_472; // @[Cat.scala 29:58]
  wire [7:0] _GEN_474 = 10'h1da == _T_7[9:0] ? 8'h0 : _GEN_473; // @[Cat.scala 29:58]
  wire [7:0] _GEN_475 = 10'h1db == _T_7[9:0] ? 8'h0 : _GEN_474; // @[Cat.scala 29:58]
  wire [7:0] _GEN_476 = 10'h1dc == _T_7[9:0] ? 8'h0 : _GEN_475; // @[Cat.scala 29:58]
  wire [7:0] _GEN_477 = 10'h1dd == _T_7[9:0] ? 8'h0 : _GEN_476; // @[Cat.scala 29:58]
  wire [7:0] _GEN_478 = 10'h1de == _T_7[9:0] ? 8'h0 : _GEN_477; // @[Cat.scala 29:58]
  wire [7:0] _GEN_479 = 10'h1df == _T_7[9:0] ? 8'h0 : _GEN_478; // @[Cat.scala 29:58]
  wire [7:0] _GEN_480 = 10'h1e0 == _T_7[9:0] ? 8'h0 : _GEN_479; // @[Cat.scala 29:58]
  wire [7:0] _GEN_481 = 10'h1e1 == _T_7[9:0] ? 8'h0 : _GEN_480; // @[Cat.scala 29:58]
  wire [7:0] _GEN_482 = 10'h1e2 == _T_7[9:0] ? 8'h0 : _GEN_481; // @[Cat.scala 29:58]
  wire [7:0] _GEN_483 = 10'h1e3 == _T_7[9:0] ? 8'h0 : _GEN_482; // @[Cat.scala 29:58]
  wire [7:0] _GEN_484 = 10'h1e4 == _T_7[9:0] ? 8'h0 : _GEN_483; // @[Cat.scala 29:58]
  wire [7:0] _GEN_485 = 10'h1e5 == _T_7[9:0] ? 8'h0 : _GEN_484; // @[Cat.scala 29:58]
  wire [7:0] _GEN_486 = 10'h1e6 == _T_7[9:0] ? 8'h0 : _GEN_485; // @[Cat.scala 29:58]
  wire [7:0] _GEN_487 = 10'h1e7 == _T_7[9:0] ? 8'h0 : _GEN_486; // @[Cat.scala 29:58]
  wire [7:0] _GEN_488 = 10'h1e8 == _T_7[9:0] ? 8'h0 : _GEN_487; // @[Cat.scala 29:58]
  wire [7:0] _GEN_489 = 10'h1e9 == _T_7[9:0] ? 8'h0 : _GEN_488; // @[Cat.scala 29:58]
  wire [7:0] _GEN_490 = 10'h1ea == _T_7[9:0] ? 8'h0 : _GEN_489; // @[Cat.scala 29:58]
  wire [7:0] _GEN_491 = 10'h1eb == _T_7[9:0] ? 8'h0 : _GEN_490; // @[Cat.scala 29:58]
  wire [7:0] _GEN_492 = 10'h1ec == _T_7[9:0] ? 8'h0 : _GEN_491; // @[Cat.scala 29:58]
  wire [7:0] _GEN_493 = 10'h1ed == _T_7[9:0] ? 8'h0 : _GEN_492; // @[Cat.scala 29:58]
  wire [7:0] _GEN_494 = 10'h1ee == _T_7[9:0] ? 8'h0 : _GEN_493; // @[Cat.scala 29:58]
  wire [7:0] _GEN_495 = 10'h1ef == _T_7[9:0] ? 8'h0 : _GEN_494; // @[Cat.scala 29:58]
  wire [7:0] _GEN_496 = 10'h1f0 == _T_7[9:0] ? 8'h0 : _GEN_495; // @[Cat.scala 29:58]
  wire [7:0] _GEN_497 = 10'h1f1 == _T_7[9:0] ? 8'h0 : _GEN_496; // @[Cat.scala 29:58]
  wire [7:0] _GEN_498 = 10'h1f2 == _T_7[9:0] ? 8'h0 : _GEN_497; // @[Cat.scala 29:58]
  wire [7:0] _GEN_499 = 10'h1f3 == _T_7[9:0] ? 8'h0 : _GEN_498; // @[Cat.scala 29:58]
  wire [7:0] _GEN_500 = 10'h1f4 == _T_7[9:0] ? 8'h0 : _GEN_499; // @[Cat.scala 29:58]
  wire [7:0] _GEN_501 = 10'h1f5 == _T_7[9:0] ? 8'h0 : _GEN_500; // @[Cat.scala 29:58]
  wire [7:0] _GEN_502 = 10'h1f6 == _T_7[9:0] ? 8'h0 : _GEN_501; // @[Cat.scala 29:58]
  wire [7:0] _GEN_503 = 10'h1f7 == _T_7[9:0] ? 8'h0 : _GEN_502; // @[Cat.scala 29:58]
  wire [7:0] _GEN_504 = 10'h1f8 == _T_7[9:0] ? 8'h0 : _GEN_503; // @[Cat.scala 29:58]
  wire [7:0] _GEN_505 = 10'h1f9 == _T_7[9:0] ? 8'h0 : _GEN_504; // @[Cat.scala 29:58]
  wire [7:0] _GEN_506 = 10'h1fa == _T_7[9:0] ? 8'h0 : _GEN_505; // @[Cat.scala 29:58]
  wire [7:0] _GEN_507 = 10'h1fb == _T_7[9:0] ? 8'h0 : _GEN_506; // @[Cat.scala 29:58]
  wire [7:0] _GEN_508 = 10'h1fc == _T_7[9:0] ? 8'h0 : _GEN_507; // @[Cat.scala 29:58]
  wire [7:0] _GEN_509 = 10'h1fd == _T_7[9:0] ? 8'h0 : _GEN_508; // @[Cat.scala 29:58]
  wire [7:0] _GEN_510 = 10'h1fe == _T_7[9:0] ? 8'h0 : _GEN_509; // @[Cat.scala 29:58]
  wire [7:0] _GEN_511 = 10'h1ff == _T_7[9:0] ? 8'h0 : _GEN_510; // @[Cat.scala 29:58]
  wire [7:0] _GEN_512 = 10'h200 == _T_7[9:0] ? 8'h0 : _GEN_511; // @[Cat.scala 29:58]
  wire [7:0] _GEN_513 = 10'h201 == _T_7[9:0] ? 8'h0 : _GEN_512; // @[Cat.scala 29:58]
  wire [7:0] _GEN_514 = 10'h202 == _T_7[9:0] ? 8'h0 : _GEN_513; // @[Cat.scala 29:58]
  wire [7:0] _GEN_515 = 10'h203 == _T_7[9:0] ? 8'h0 : _GEN_514; // @[Cat.scala 29:58]
  wire [7:0] _GEN_516 = 10'h204 == _T_7[9:0] ? 8'h0 : _GEN_515; // @[Cat.scala 29:58]
  wire [7:0] _GEN_517 = 10'h205 == _T_7[9:0] ? 8'h0 : _GEN_516; // @[Cat.scala 29:58]
  wire [7:0] _GEN_518 = 10'h206 == _T_7[9:0] ? 8'h0 : _GEN_517; // @[Cat.scala 29:58]
  wire [7:0] _GEN_519 = 10'h207 == _T_7[9:0] ? 8'h0 : _GEN_518; // @[Cat.scala 29:58]
  wire [7:0] _GEN_520 = 10'h208 == _T_7[9:0] ? 8'h0 : _GEN_519; // @[Cat.scala 29:58]
  wire [7:0] _GEN_521 = 10'h209 == _T_7[9:0] ? 8'h0 : _GEN_520; // @[Cat.scala 29:58]
  wire [7:0] _GEN_522 = 10'h20a == _T_7[9:0] ? 8'h0 : _GEN_521; // @[Cat.scala 29:58]
  wire [7:0] _GEN_523 = 10'h20b == _T_7[9:0] ? 8'h0 : _GEN_522; // @[Cat.scala 29:58]
  wire [7:0] _GEN_525 = 10'h1 == pc[9:0] ? 8'h21 : 8'h97; // @[Cat.scala 29:58]
  wire [7:0] _GEN_526 = 10'h2 == pc[9:0] ? 8'h0 : _GEN_525; // @[Cat.scala 29:58]
  wire [7:0] _GEN_527 = 10'h3 == pc[9:0] ? 8'h0 : _GEN_526; // @[Cat.scala 29:58]
  wire [7:0] _GEN_528 = 10'h4 == pc[9:0] ? 8'h93 : _GEN_527; // @[Cat.scala 29:58]
  wire [7:0] _GEN_529 = 10'h5 == pc[9:0] ? 8'h81 : _GEN_528; // @[Cat.scala 29:58]
  wire [7:0] _GEN_530 = 10'h6 == pc[9:0] ? 8'h1 : _GEN_529; // @[Cat.scala 29:58]
  wire [7:0] _GEN_531 = 10'h7 == pc[9:0] ? 8'h97 : _GEN_530; // @[Cat.scala 29:58]
  wire [7:0] _GEN_532 = 10'h8 == pc[9:0] ? 8'h17 : _GEN_531; // @[Cat.scala 29:58]
  wire [7:0] _GEN_533 = 10'h9 == pc[9:0] ? 8'h11 : _GEN_532; // @[Cat.scala 29:58]
  wire [7:0] _GEN_534 = 10'ha == pc[9:0] ? 8'h0 : _GEN_533; // @[Cat.scala 29:58]
  wire [7:0] _GEN_535 = 10'hb == pc[9:0] ? 8'h0 : _GEN_534; // @[Cat.scala 29:58]
  wire [7:0] _GEN_536 = 10'hc == pc[9:0] ? 8'h13 : _GEN_535; // @[Cat.scala 29:58]
  wire [7:0] _GEN_537 = 10'hd == pc[9:0] ? 8'h1 : _GEN_536; // @[Cat.scala 29:58]
  wire [7:0] _GEN_538 = 10'he == pc[9:0] ? 8'h81 : _GEN_537; // @[Cat.scala 29:58]
  wire [7:0] _GEN_539 = 10'hf == pc[9:0] ? 8'hff : _GEN_538; // @[Cat.scala 29:58]
  wire [7:0] _GEN_540 = 10'h10 == pc[9:0] ? 8'h33 : _GEN_539; // @[Cat.scala 29:58]
  wire [7:0] _GEN_541 = 10'h11 == pc[9:0] ? 8'h4 : _GEN_540; // @[Cat.scala 29:58]
  wire [7:0] _GEN_542 = 10'h12 == pc[9:0] ? 8'h1 : _GEN_541; // @[Cat.scala 29:58]
  wire [7:0] _GEN_543 = 10'h13 == pc[9:0] ? 8'h0 : _GEN_542; // @[Cat.scala 29:58]
  wire [7:0] _GEN_544 = 10'h14 == pc[9:0] ? 8'h6f : _GEN_543; // @[Cat.scala 29:58]
  wire [7:0] _GEN_545 = 10'h15 == pc[9:0] ? 8'h0 : _GEN_544; // @[Cat.scala 29:58]
  wire [7:0] _GEN_546 = 10'h16 == pc[9:0] ? 8'h80 : _GEN_545; // @[Cat.scala 29:58]
  wire [7:0] _GEN_547 = 10'h17 == pc[9:0] ? 8'h9 : _GEN_546; // @[Cat.scala 29:58]
  wire [7:0] _GEN_548 = 10'h18 == pc[9:0] ? 8'h13 : _GEN_547; // @[Cat.scala 29:58]
  wire [7:0] _GEN_549 = 10'h19 == pc[9:0] ? 8'h1 : _GEN_548; // @[Cat.scala 29:58]
  wire [7:0] _GEN_550 = 10'h1a == pc[9:0] ? 8'h1 : _GEN_549; // @[Cat.scala 29:58]
  wire [7:0] _GEN_551 = 10'h1b == pc[9:0] ? 8'hfe : _GEN_550; // @[Cat.scala 29:58]
  wire [7:0] _GEN_552 = 10'h1c == pc[9:0] ? 8'h23 : _GEN_551; // @[Cat.scala 29:58]
  wire [7:0] _GEN_553 = 10'h1d == pc[9:0] ? 8'h2e : _GEN_552; // @[Cat.scala 29:58]
  wire [7:0] _GEN_554 = 10'h1e == pc[9:0] ? 8'h81 : _GEN_553; // @[Cat.scala 29:58]
  wire [7:0] _GEN_555 = 10'h1f == pc[9:0] ? 8'h0 : _GEN_554; // @[Cat.scala 29:58]
  wire [7:0] _GEN_556 = 10'h20 == pc[9:0] ? 8'h13 : _GEN_555; // @[Cat.scala 29:58]
  wire [7:0] _GEN_557 = 10'h21 == pc[9:0] ? 8'h4 : _GEN_556; // @[Cat.scala 29:58]
  wire [7:0] _GEN_558 = 10'h22 == pc[9:0] ? 8'h1 : _GEN_557; // @[Cat.scala 29:58]
  wire [7:0] _GEN_559 = 10'h23 == pc[9:0] ? 8'h2 : _GEN_558; // @[Cat.scala 29:58]
  wire [7:0] _GEN_560 = 10'h24 == pc[9:0] ? 8'hb7 : _GEN_559; // @[Cat.scala 29:58]
  wire [7:0] _GEN_561 = 10'h25 == pc[9:0] ? 8'h27 : _GEN_560; // @[Cat.scala 29:58]
  wire [7:0] _GEN_562 = 10'h26 == pc[9:0] ? 8'h0 : _GEN_561; // @[Cat.scala 29:58]
  wire [7:0] _GEN_563 = 10'h27 == pc[9:0] ? 8'h0 : _GEN_562; // @[Cat.scala 29:58]
  wire [7:0] _GEN_564 = 10'h28 == pc[9:0] ? 8'h93 : _GEN_563; // @[Cat.scala 29:58]
  wire [7:0] _GEN_565 = 10'h29 == pc[9:0] ? 8'h87 : _GEN_564; // @[Cat.scala 29:58]
  wire [7:0] _GEN_566 = 10'h2a == pc[9:0] ? 8'h7 : _GEN_565; // @[Cat.scala 29:58]
  wire [7:0] _GEN_567 = 10'h2b == pc[9:0] ? 8'h20 : _GEN_566; // @[Cat.scala 29:58]
  wire [7:0] _GEN_568 = 10'h2c == pc[9:0] ? 8'h23 : _GEN_567; // @[Cat.scala 29:58]
  wire [7:0] _GEN_569 = 10'h2d == pc[9:0] ? 8'h26 : _GEN_568; // @[Cat.scala 29:58]
  wire [7:0] _GEN_570 = 10'h2e == pc[9:0] ? 8'hf4 : _GEN_569; // @[Cat.scala 29:58]
  wire [7:0] _GEN_571 = 10'h2f == pc[9:0] ? 8'hfe : _GEN_570; // @[Cat.scala 29:58]
  wire [7:0] _GEN_572 = 10'h30 == pc[9:0] ? 8'h83 : _GEN_571; // @[Cat.scala 29:58]
  wire [7:0] _GEN_573 = 10'h31 == pc[9:0] ? 8'h27 : _GEN_572; // @[Cat.scala 29:58]
  wire [7:0] _GEN_574 = 10'h32 == pc[9:0] ? 8'hc4 : _GEN_573; // @[Cat.scala 29:58]
  wire [7:0] _GEN_575 = 10'h33 == pc[9:0] ? 8'hfe : _GEN_574; // @[Cat.scala 29:58]
  wire [7:0] _GEN_576 = 10'h34 == pc[9:0] ? 8'h83 : _GEN_575; // @[Cat.scala 29:58]
  wire [7:0] _GEN_577 = 10'h35 == pc[9:0] ? 8'ha7 : _GEN_576; // @[Cat.scala 29:58]
  wire [7:0] _GEN_578 = 10'h36 == pc[9:0] ? 8'h7 : _GEN_577; // @[Cat.scala 29:58]
  wire [7:0] _GEN_579 = 10'h37 == pc[9:0] ? 8'h0 : _GEN_578; // @[Cat.scala 29:58]
  wire [7:0] _GEN_580 = 10'h38 == pc[9:0] ? 8'h13 : _GEN_579; // @[Cat.scala 29:58]
  wire [7:0] _GEN_581 = 10'h39 == pc[9:0] ? 8'h85 : _GEN_580; // @[Cat.scala 29:58]
  wire [7:0] _GEN_582 = 10'h3a == pc[9:0] ? 8'h7 : _GEN_581; // @[Cat.scala 29:58]
  wire [7:0] _GEN_583 = 10'h3b == pc[9:0] ? 8'h0 : _GEN_582; // @[Cat.scala 29:58]
  wire [7:0] _GEN_584 = 10'h3c == pc[9:0] ? 8'h3 : _GEN_583; // @[Cat.scala 29:58]
  wire [7:0] _GEN_585 = 10'h3d == pc[9:0] ? 8'h24 : _GEN_584; // @[Cat.scala 29:58]
  wire [7:0] _GEN_586 = 10'h3e == pc[9:0] ? 8'hc1 : _GEN_585; // @[Cat.scala 29:58]
  wire [7:0] _GEN_587 = 10'h3f == pc[9:0] ? 8'h1 : _GEN_586; // @[Cat.scala 29:58]
  wire [7:0] _GEN_588 = 10'h40 == pc[9:0] ? 8'h13 : _GEN_587; // @[Cat.scala 29:58]
  wire [7:0] _GEN_589 = 10'h41 == pc[9:0] ? 8'h1 : _GEN_588; // @[Cat.scala 29:58]
  wire [7:0] _GEN_590 = 10'h42 == pc[9:0] ? 8'h1 : _GEN_589; // @[Cat.scala 29:58]
  wire [7:0] _GEN_591 = 10'h43 == pc[9:0] ? 8'h2 : _GEN_590; // @[Cat.scala 29:58]
  wire [7:0] _GEN_592 = 10'h44 == pc[9:0] ? 8'h67 : _GEN_591; // @[Cat.scala 29:58]
  wire [7:0] _GEN_593 = 10'h45 == pc[9:0] ? 8'h80 : _GEN_592; // @[Cat.scala 29:58]
  wire [7:0] _GEN_594 = 10'h46 == pc[9:0] ? 8'h0 : _GEN_593; // @[Cat.scala 29:58]
  wire [7:0] _GEN_595 = 10'h47 == pc[9:0] ? 8'h0 : _GEN_594; // @[Cat.scala 29:58]
  wire [7:0] _GEN_596 = 10'h48 == pc[9:0] ? 8'h13 : _GEN_595; // @[Cat.scala 29:58]
  wire [7:0] _GEN_597 = 10'h49 == pc[9:0] ? 8'h1 : _GEN_596; // @[Cat.scala 29:58]
  wire [7:0] _GEN_598 = 10'h4a == pc[9:0] ? 8'h1 : _GEN_597; // @[Cat.scala 29:58]
  wire [7:0] _GEN_599 = 10'h4b == pc[9:0] ? 8'hfe : _GEN_598; // @[Cat.scala 29:58]
  wire [7:0] _GEN_600 = 10'h4c == pc[9:0] ? 8'h23 : _GEN_599; // @[Cat.scala 29:58]
  wire [7:0] _GEN_601 = 10'h4d == pc[9:0] ? 8'h2e : _GEN_600; // @[Cat.scala 29:58]
  wire [7:0] _GEN_602 = 10'h4e == pc[9:0] ? 8'h81 : _GEN_601; // @[Cat.scala 29:58]
  wire [7:0] _GEN_603 = 10'h4f == pc[9:0] ? 8'h0 : _GEN_602; // @[Cat.scala 29:58]
  wire [7:0] _GEN_604 = 10'h50 == pc[9:0] ? 8'h13 : _GEN_603; // @[Cat.scala 29:58]
  wire [7:0] _GEN_605 = 10'h51 == pc[9:0] ? 8'h4 : _GEN_604; // @[Cat.scala 29:58]
  wire [7:0] _GEN_606 = 10'h52 == pc[9:0] ? 8'h1 : _GEN_605; // @[Cat.scala 29:58]
  wire [7:0] _GEN_607 = 10'h53 == pc[9:0] ? 8'h2 : _GEN_606; // @[Cat.scala 29:58]
  wire [7:0] _GEN_608 = 10'h54 == pc[9:0] ? 8'hb7 : _GEN_607; // @[Cat.scala 29:58]
  wire [7:0] _GEN_609 = 10'h55 == pc[9:0] ? 8'h27 : _GEN_608; // @[Cat.scala 29:58]
  wire [7:0] _GEN_610 = 10'h56 == pc[9:0] ? 8'h0 : _GEN_609; // @[Cat.scala 29:58]
  wire [7:0] _GEN_611 = 10'h57 == pc[9:0] ? 8'h0 : _GEN_610; // @[Cat.scala 29:58]
  wire [7:0] _GEN_612 = 10'h58 == pc[9:0] ? 8'h93 : _GEN_611; // @[Cat.scala 29:58]
  wire [7:0] _GEN_613 = 10'h59 == pc[9:0] ? 8'h87 : _GEN_612; // @[Cat.scala 29:58]
  wire [7:0] _GEN_614 = 10'h5a == pc[9:0] ? 8'h7 : _GEN_613; // @[Cat.scala 29:58]
  wire [7:0] _GEN_615 = 10'h5b == pc[9:0] ? 8'h10 : _GEN_614; // @[Cat.scala 29:58]
  wire [7:0] _GEN_616 = 10'h5c == pc[9:0] ? 8'h23 : _GEN_615; // @[Cat.scala 29:58]
  wire [7:0] _GEN_617 = 10'h5d == pc[9:0] ? 8'h26 : _GEN_616; // @[Cat.scala 29:58]
  wire [7:0] _GEN_618 = 10'h5e == pc[9:0] ? 8'hf4 : _GEN_617; // @[Cat.scala 29:58]
  wire [7:0] _GEN_619 = 10'h5f == pc[9:0] ? 8'hfe : _GEN_618; // @[Cat.scala 29:58]
  wire [7:0] _GEN_620 = 10'h60 == pc[9:0] ? 8'h83 : _GEN_619; // @[Cat.scala 29:58]
  wire [7:0] _GEN_621 = 10'h61 == pc[9:0] ? 8'h27 : _GEN_620; // @[Cat.scala 29:58]
  wire [7:0] _GEN_622 = 10'h62 == pc[9:0] ? 8'hc4 : _GEN_621; // @[Cat.scala 29:58]
  wire [7:0] _GEN_623 = 10'h63 == pc[9:0] ? 8'hfe : _GEN_622; // @[Cat.scala 29:58]
  wire [7:0] _GEN_624 = 10'h64 == pc[9:0] ? 8'h83 : _GEN_623; // @[Cat.scala 29:58]
  wire [7:0] _GEN_625 = 10'h65 == pc[9:0] ? 8'ha7 : _GEN_624; // @[Cat.scala 29:58]
  wire [7:0] _GEN_626 = 10'h66 == pc[9:0] ? 8'h7 : _GEN_625; // @[Cat.scala 29:58]
  wire [7:0] _GEN_627 = 10'h67 == pc[9:0] ? 8'h0 : _GEN_626; // @[Cat.scala 29:58]
  wire [7:0] _GEN_628 = 10'h68 == pc[9:0] ? 8'h13 : _GEN_627; // @[Cat.scala 29:58]
  wire [7:0] _GEN_629 = 10'h69 == pc[9:0] ? 8'h85 : _GEN_628; // @[Cat.scala 29:58]
  wire [7:0] _GEN_630 = 10'h6a == pc[9:0] ? 8'h7 : _GEN_629; // @[Cat.scala 29:58]
  wire [7:0] _GEN_631 = 10'h6b == pc[9:0] ? 8'h0 : _GEN_630; // @[Cat.scala 29:58]
  wire [7:0] _GEN_632 = 10'h6c == pc[9:0] ? 8'h3 : _GEN_631; // @[Cat.scala 29:58]
  wire [7:0] _GEN_633 = 10'h6d == pc[9:0] ? 8'h24 : _GEN_632; // @[Cat.scala 29:58]
  wire [7:0] _GEN_634 = 10'h6e == pc[9:0] ? 8'hc1 : _GEN_633; // @[Cat.scala 29:58]
  wire [7:0] _GEN_635 = 10'h6f == pc[9:0] ? 8'h1 : _GEN_634; // @[Cat.scala 29:58]
  wire [7:0] _GEN_636 = 10'h70 == pc[9:0] ? 8'h13 : _GEN_635; // @[Cat.scala 29:58]
  wire [7:0] _GEN_637 = 10'h71 == pc[9:0] ? 8'h1 : _GEN_636; // @[Cat.scala 29:58]
  wire [7:0] _GEN_638 = 10'h72 == pc[9:0] ? 8'h1 : _GEN_637; // @[Cat.scala 29:58]
  wire [7:0] _GEN_639 = 10'h73 == pc[9:0] ? 8'h2 : _GEN_638; // @[Cat.scala 29:58]
  wire [7:0] _GEN_640 = 10'h74 == pc[9:0] ? 8'h67 : _GEN_639; // @[Cat.scala 29:58]
  wire [7:0] _GEN_641 = 10'h75 == pc[9:0] ? 8'h80 : _GEN_640; // @[Cat.scala 29:58]
  wire [7:0] _GEN_642 = 10'h76 == pc[9:0] ? 8'h0 : _GEN_641; // @[Cat.scala 29:58]
  wire [7:0] _GEN_643 = 10'h77 == pc[9:0] ? 8'h0 : _GEN_642; // @[Cat.scala 29:58]
  wire [7:0] _GEN_644 = 10'h78 == pc[9:0] ? 8'h13 : _GEN_643; // @[Cat.scala 29:58]
  wire [7:0] _GEN_645 = 10'h79 == pc[9:0] ? 8'h1 : _GEN_644; // @[Cat.scala 29:58]
  wire [7:0] _GEN_646 = 10'h7a == pc[9:0] ? 8'h1 : _GEN_645; // @[Cat.scala 29:58]
  wire [7:0] _GEN_647 = 10'h7b == pc[9:0] ? 8'hfd : _GEN_646; // @[Cat.scala 29:58]
  wire [7:0] _GEN_648 = 10'h7c == pc[9:0] ? 8'h23 : _GEN_647; // @[Cat.scala 29:58]
  wire [7:0] _GEN_649 = 10'h7d == pc[9:0] ? 8'h26 : _GEN_648; // @[Cat.scala 29:58]
  wire [7:0] _GEN_650 = 10'h7e == pc[9:0] ? 8'h81 : _GEN_649; // @[Cat.scala 29:58]
  wire [7:0] _GEN_651 = 10'h7f == pc[9:0] ? 8'h2 : _GEN_650; // @[Cat.scala 29:58]
  wire [7:0] _GEN_652 = 10'h80 == pc[9:0] ? 8'h13 : _GEN_651; // @[Cat.scala 29:58]
  wire [7:0] _GEN_653 = 10'h81 == pc[9:0] ? 8'h4 : _GEN_652; // @[Cat.scala 29:58]
  wire [7:0] _GEN_654 = 10'h82 == pc[9:0] ? 8'h1 : _GEN_653; // @[Cat.scala 29:58]
  wire [7:0] _GEN_655 = 10'h83 == pc[9:0] ? 8'h3 : _GEN_654; // @[Cat.scala 29:58]
  wire [7:0] _GEN_656 = 10'h84 == pc[9:0] ? 8'h23 : _GEN_655; // @[Cat.scala 29:58]
  wire [7:0] _GEN_657 = 10'h85 == pc[9:0] ? 8'h2e : _GEN_656; // @[Cat.scala 29:58]
  wire [7:0] _GEN_658 = 10'h86 == pc[9:0] ? 8'ha4 : _GEN_657; // @[Cat.scala 29:58]
  wire [7:0] _GEN_659 = 10'h87 == pc[9:0] ? 8'hfc : _GEN_658; // @[Cat.scala 29:58]
  wire [7:0] _GEN_660 = 10'h88 == pc[9:0] ? 8'hb7 : _GEN_659; // @[Cat.scala 29:58]
  wire [7:0] _GEN_661 = 10'h89 == pc[9:0] ? 8'h27 : _GEN_660; // @[Cat.scala 29:58]
  wire [7:0] _GEN_662 = 10'h8a == pc[9:0] ? 8'h0 : _GEN_661; // @[Cat.scala 29:58]
  wire [7:0] _GEN_663 = 10'h8b == pc[9:0] ? 8'h0 : _GEN_662; // @[Cat.scala 29:58]
  wire [7:0] _GEN_664 = 10'h8c == pc[9:0] ? 8'h23 : _GEN_663; // @[Cat.scala 29:58]
  wire [7:0] _GEN_665 = 10'h8d == pc[9:0] ? 8'h26 : _GEN_664; // @[Cat.scala 29:58]
  wire [7:0] _GEN_666 = 10'h8e == pc[9:0] ? 8'hf4 : _GEN_665; // @[Cat.scala 29:58]
  wire [7:0] _GEN_667 = 10'h8f == pc[9:0] ? 8'hfe : _GEN_666; // @[Cat.scala 29:58]
  wire [7:0] _GEN_668 = 10'h90 == pc[9:0] ? 8'h83 : _GEN_667; // @[Cat.scala 29:58]
  wire [7:0] _GEN_669 = 10'h91 == pc[9:0] ? 8'h27 : _GEN_668; // @[Cat.scala 29:58]
  wire [7:0] _GEN_670 = 10'h92 == pc[9:0] ? 8'hc4 : _GEN_669; // @[Cat.scala 29:58]
  wire [7:0] _GEN_671 = 10'h93 == pc[9:0] ? 8'hfe : _GEN_670; // @[Cat.scala 29:58]
  wire [7:0] _GEN_672 = 10'h94 == pc[9:0] ? 8'h3 : _GEN_671; // @[Cat.scala 29:58]
  wire [7:0] _GEN_673 = 10'h95 == pc[9:0] ? 8'h27 : _GEN_672; // @[Cat.scala 29:58]
  wire [7:0] _GEN_674 = 10'h96 == pc[9:0] ? 8'hc4 : _GEN_673; // @[Cat.scala 29:58]
  wire [7:0] _GEN_675 = 10'h97 == pc[9:0] ? 8'hfd : _GEN_674; // @[Cat.scala 29:58]
  wire [7:0] _GEN_676 = 10'h98 == pc[9:0] ? 8'h23 : _GEN_675; // @[Cat.scala 29:58]
  wire [7:0] _GEN_677 = 10'h99 == pc[9:0] ? 8'ha0 : _GEN_676; // @[Cat.scala 29:58]
  wire [7:0] _GEN_678 = 10'h9a == pc[9:0] ? 8'he7 : _GEN_677; // @[Cat.scala 29:58]
  wire [7:0] _GEN_679 = 10'h9b == pc[9:0] ? 8'h0 : _GEN_678; // @[Cat.scala 29:58]
  wire [7:0] _GEN_680 = 10'h9c == pc[9:0] ? 8'h13 : _GEN_679; // @[Cat.scala 29:58]
  wire [7:0] _GEN_681 = 10'h9d == pc[9:0] ? 8'h0 : _GEN_680; // @[Cat.scala 29:58]
  wire [7:0] _GEN_682 = 10'h9e == pc[9:0] ? 8'h0 : _GEN_681; // @[Cat.scala 29:58]
  wire [7:0] _GEN_683 = 10'h9f == pc[9:0] ? 8'h0 : _GEN_682; // @[Cat.scala 29:58]
  wire [7:0] _GEN_684 = 10'ha0 == pc[9:0] ? 8'h3 : _GEN_683; // @[Cat.scala 29:58]
  wire [7:0] _GEN_685 = 10'ha1 == pc[9:0] ? 8'h24 : _GEN_684; // @[Cat.scala 29:58]
  wire [7:0] _GEN_686 = 10'ha2 == pc[9:0] ? 8'hc1 : _GEN_685; // @[Cat.scala 29:58]
  wire [7:0] _GEN_687 = 10'ha3 == pc[9:0] ? 8'h2 : _GEN_686; // @[Cat.scala 29:58]
  wire [7:0] _GEN_688 = 10'ha4 == pc[9:0] ? 8'h13 : _GEN_687; // @[Cat.scala 29:58]
  wire [7:0] _GEN_689 = 10'ha5 == pc[9:0] ? 8'h1 : _GEN_688; // @[Cat.scala 29:58]
  wire [7:0] _GEN_690 = 10'ha6 == pc[9:0] ? 8'h1 : _GEN_689; // @[Cat.scala 29:58]
  wire [7:0] _GEN_691 = 10'ha7 == pc[9:0] ? 8'h3 : _GEN_690; // @[Cat.scala 29:58]
  wire [7:0] _GEN_692 = 10'ha8 == pc[9:0] ? 8'h67 : _GEN_691; // @[Cat.scala 29:58]
  wire [7:0] _GEN_693 = 10'ha9 == pc[9:0] ? 8'h80 : _GEN_692; // @[Cat.scala 29:58]
  wire [7:0] _GEN_694 = 10'haa == pc[9:0] ? 8'h0 : _GEN_693; // @[Cat.scala 29:58]
  wire [7:0] _GEN_695 = 10'hab == pc[9:0] ? 8'h0 : _GEN_694; // @[Cat.scala 29:58]
  wire [7:0] _GEN_696 = 10'hac == pc[9:0] ? 8'h13 : _GEN_695; // @[Cat.scala 29:58]
  wire [7:0] _GEN_697 = 10'had == pc[9:0] ? 8'h1 : _GEN_696; // @[Cat.scala 29:58]
  wire [7:0] _GEN_698 = 10'hae == pc[9:0] ? 8'h1 : _GEN_697; // @[Cat.scala 29:58]
  wire [7:0] _GEN_699 = 10'haf == pc[9:0] ? 8'hfe : _GEN_698; // @[Cat.scala 29:58]
  wire [7:0] _GEN_700 = 10'hb0 == pc[9:0] ? 8'h23 : _GEN_699; // @[Cat.scala 29:58]
  wire [7:0] _GEN_701 = 10'hb1 == pc[9:0] ? 8'h2e : _GEN_700; // @[Cat.scala 29:58]
  wire [7:0] _GEN_702 = 10'hb2 == pc[9:0] ? 8'h11 : _GEN_701; // @[Cat.scala 29:58]
  wire [7:0] _GEN_703 = 10'hb3 == pc[9:0] ? 8'h0 : _GEN_702; // @[Cat.scala 29:58]
  wire [7:0] _GEN_704 = 10'hb4 == pc[9:0] ? 8'h23 : _GEN_703; // @[Cat.scala 29:58]
  wire [7:0] _GEN_705 = 10'hb5 == pc[9:0] ? 8'h2c : _GEN_704; // @[Cat.scala 29:58]
  wire [7:0] _GEN_706 = 10'hb6 == pc[9:0] ? 8'h81 : _GEN_705; // @[Cat.scala 29:58]
  wire [7:0] _GEN_707 = 10'hb7 == pc[9:0] ? 8'h0 : _GEN_706; // @[Cat.scala 29:58]
  wire [7:0] _GEN_708 = 10'hb8 == pc[9:0] ? 8'h13 : _GEN_707; // @[Cat.scala 29:58]
  wire [7:0] _GEN_709 = 10'hb9 == pc[9:0] ? 8'h4 : _GEN_708; // @[Cat.scala 29:58]
  wire [7:0] _GEN_710 = 10'hba == pc[9:0] ? 8'h1 : _GEN_709; // @[Cat.scala 29:58]
  wire [7:0] _GEN_711 = 10'hbb == pc[9:0] ? 8'h2 : _GEN_710; // @[Cat.scala 29:58]
  wire [7:0] _GEN_712 = 10'hbc == pc[9:0] ? 8'h23 : _GEN_711; // @[Cat.scala 29:58]
  wire [7:0] _GEN_713 = 10'hbd == pc[9:0] ? 8'h26 : _GEN_712; // @[Cat.scala 29:58]
  wire [7:0] _GEN_714 = 10'hbe == pc[9:0] ? 8'h4 : _GEN_713; // @[Cat.scala 29:58]
  wire [7:0] _GEN_715 = 10'hbf == pc[9:0] ? 8'hfe : _GEN_714; // @[Cat.scala 29:58]
  wire [7:0] _GEN_716 = 10'hc0 == pc[9:0] ? 8'hb7 : _GEN_715; // @[Cat.scala 29:58]
  wire [7:0] _GEN_717 = 10'hc1 == pc[9:0] ? 8'hc7 : _GEN_716; // @[Cat.scala 29:58]
  wire [7:0] _GEN_718 = 10'hc2 == pc[9:0] ? 8'h0 : _GEN_717; // @[Cat.scala 29:58]
  wire [7:0] _GEN_719 = 10'hc3 == pc[9:0] ? 8'h0 : _GEN_718; // @[Cat.scala 29:58]
  wire [7:0] _GEN_720 = 10'hc4 == pc[9:0] ? 8'h13 : _GEN_719; // @[Cat.scala 29:58]
  wire [7:0] _GEN_721 = 10'hc5 == pc[9:0] ? 8'h85 : _GEN_720; // @[Cat.scala 29:58]
  wire [7:0] _GEN_722 = 10'hc6 == pc[9:0] ? 8'hf7 : _GEN_721; // @[Cat.scala 29:58]
  wire [7:0] _GEN_723 = 10'hc7 == pc[9:0] ? 8'hee : _GEN_722; // @[Cat.scala 29:58]
  wire [7:0] _GEN_724 = 10'hc8 == pc[9:0] ? 8'hef : _GEN_723; // @[Cat.scala 29:58]
  wire [7:0] _GEN_725 = 10'hc9 == pc[9:0] ? 8'hf0 : _GEN_724; // @[Cat.scala 29:58]
  wire [7:0] _GEN_726 = 10'hca == pc[9:0] ? 8'h1f : _GEN_725; // @[Cat.scala 29:58]
  wire [7:0] _GEN_727 = 10'hcb == pc[9:0] ? 8'hfb : _GEN_726; // @[Cat.scala 29:58]
  wire [7:0] _GEN_728 = 10'hcc == pc[9:0] ? 8'h23 : _GEN_727; // @[Cat.scala 29:58]
  wire [7:0] _GEN_729 = 10'hcd == pc[9:0] ? 8'h26 : _GEN_728; // @[Cat.scala 29:58]
  wire [7:0] _GEN_730 = 10'hce == pc[9:0] ? 8'h4 : _GEN_729; // @[Cat.scala 29:58]
  wire [7:0] _GEN_731 = 10'hcf == pc[9:0] ? 8'hfe : _GEN_730; // @[Cat.scala 29:58]
  wire [7:0] _GEN_732 = 10'hd0 == pc[9:0] ? 8'h6f : _GEN_731; // @[Cat.scala 29:58]
  wire [7:0] _GEN_733 = 10'hd1 == pc[9:0] ? 8'h0 : _GEN_732; // @[Cat.scala 29:58]
  wire [7:0] _GEN_734 = 10'hd2 == pc[9:0] ? 8'h0 : _GEN_733; // @[Cat.scala 29:58]
  wire [7:0] _GEN_735 = 10'hd3 == pc[9:0] ? 8'h1 : _GEN_734; // @[Cat.scala 29:58]
  wire [7:0] _GEN_736 = 10'hd4 == pc[9:0] ? 8'h83 : _GEN_735; // @[Cat.scala 29:58]
  wire [7:0] _GEN_737 = 10'hd5 == pc[9:0] ? 8'h27 : _GEN_736; // @[Cat.scala 29:58]
  wire [7:0] _GEN_738 = 10'hd6 == pc[9:0] ? 8'hc4 : _GEN_737; // @[Cat.scala 29:58]
  wire [7:0] _GEN_739 = 10'hd7 == pc[9:0] ? 8'hfe : _GEN_738; // @[Cat.scala 29:58]
  wire [7:0] _GEN_740 = 10'hd8 == pc[9:0] ? 8'h93 : _GEN_739; // @[Cat.scala 29:58]
  wire [7:0] _GEN_741 = 10'hd9 == pc[9:0] ? 8'h87 : _GEN_740; // @[Cat.scala 29:58]
  wire [7:0] _GEN_742 = 10'hda == pc[9:0] ? 8'h17 : _GEN_741; // @[Cat.scala 29:58]
  wire [7:0] _GEN_743 = 10'hdb == pc[9:0] ? 8'h0 : _GEN_742; // @[Cat.scala 29:58]
  wire [7:0] _GEN_744 = 10'hdc == pc[9:0] ? 8'h23 : _GEN_743; // @[Cat.scala 29:58]
  wire [7:0] _GEN_745 = 10'hdd == pc[9:0] ? 8'h26 : _GEN_744; // @[Cat.scala 29:58]
  wire [7:0] _GEN_746 = 10'hde == pc[9:0] ? 8'hf4 : _GEN_745; // @[Cat.scala 29:58]
  wire [7:0] _GEN_747 = 10'hdf == pc[9:0] ? 8'hfe : _GEN_746; // @[Cat.scala 29:58]
  wire [7:0] _GEN_748 = 10'he0 == pc[9:0] ? 8'h3 : _GEN_747; // @[Cat.scala 29:58]
  wire [7:0] _GEN_749 = 10'he1 == pc[9:0] ? 8'h27 : _GEN_748; // @[Cat.scala 29:58]
  wire [7:0] _GEN_750 = 10'he2 == pc[9:0] ? 8'hc4 : _GEN_749; // @[Cat.scala 29:58]
  wire [7:0] _GEN_751 = 10'he3 == pc[9:0] ? 8'hfe : _GEN_750; // @[Cat.scala 29:58]
  wire [7:0] _GEN_752 = 10'he4 == pc[9:0] ? 8'hb7 : _GEN_751; // @[Cat.scala 29:58]
  wire [7:0] _GEN_753 = 10'he5 == pc[9:0] ? 8'h17 : _GEN_752; // @[Cat.scala 29:58]
  wire [7:0] _GEN_754 = 10'he6 == pc[9:0] ? 8'h7a : _GEN_753; // @[Cat.scala 29:58]
  wire [7:0] _GEN_755 = 10'he7 == pc[9:0] ? 8'h0 : _GEN_754; // @[Cat.scala 29:58]
  wire [7:0] _GEN_756 = 10'he8 == pc[9:0] ? 8'h93 : _GEN_755; // @[Cat.scala 29:58]
  wire [7:0] _GEN_757 = 10'he9 == pc[9:0] ? 8'h87 : _GEN_756; // @[Cat.scala 29:58]
  wire [7:0] _GEN_758 = 10'hea == pc[9:0] ? 8'hf7 : _GEN_757; // @[Cat.scala 29:58]
  wire [7:0] _GEN_759 = 10'heb == pc[9:0] ? 8'h1f : _GEN_758; // @[Cat.scala 29:58]
  wire [7:0] _GEN_760 = 10'hec == pc[9:0] ? 8'he3 : _GEN_759; // @[Cat.scala 29:58]
  wire [7:0] _GEN_761 = 10'hed == pc[9:0] ? 8'hd4 : _GEN_760; // @[Cat.scala 29:58]
  wire [7:0] _GEN_762 = 10'hee == pc[9:0] ? 8'he7 : _GEN_761; // @[Cat.scala 29:58]
  wire [7:0] _GEN_763 = 10'hef == pc[9:0] ? 8'hfe : _GEN_762; // @[Cat.scala 29:58]
  wire [7:0] _GEN_764 = 10'hf0 == pc[9:0] ? 8'h13 : _GEN_763; // @[Cat.scala 29:58]
  wire [7:0] _GEN_765 = 10'hf1 == pc[9:0] ? 8'h5 : _GEN_764; // @[Cat.scala 29:58]
  wire [7:0] _GEN_766 = 10'hf2 == pc[9:0] ? 8'h0 : _GEN_765; // @[Cat.scala 29:58]
  wire [7:0] _GEN_767 = 10'hf3 == pc[9:0] ? 8'h0 : _GEN_766; // @[Cat.scala 29:58]
  wire [7:0] _GEN_768 = 10'hf4 == pc[9:0] ? 8'hef : _GEN_767; // @[Cat.scala 29:58]
  wire [7:0] _GEN_769 = 10'hf5 == pc[9:0] ? 8'hf0 : _GEN_768; // @[Cat.scala 29:58]
  wire [7:0] _GEN_770 = 10'hf6 == pc[9:0] ? 8'h5f : _GEN_769; // @[Cat.scala 29:58]
  wire [7:0] _GEN_771 = 10'hf7 == pc[9:0] ? 8'hf8 : _GEN_770; // @[Cat.scala 29:58]
  wire [7:0] _GEN_772 = 10'hf8 == pc[9:0] ? 8'hef : _GEN_771; // @[Cat.scala 29:58]
  wire [7:0] _GEN_773 = 10'hf9 == pc[9:0] ? 8'hf0 : _GEN_772; // @[Cat.scala 29:58]
  wire [7:0] _GEN_774 = 10'hfa == pc[9:0] ? 8'h1f : _GEN_773; // @[Cat.scala 29:58]
  wire [7:0] _GEN_775 = 10'hfb == pc[9:0] ? 8'hf5 : _GEN_774; // @[Cat.scala 29:58]
  wire [7:0] _GEN_776 = 10'hfc == pc[9:0] ? 8'h93 : _GEN_775; // @[Cat.scala 29:58]
  wire [7:0] _GEN_777 = 10'hfd == pc[9:0] ? 8'h7 : _GEN_776; // @[Cat.scala 29:58]
  wire [7:0] _GEN_778 = 10'hfe == pc[9:0] ? 8'h5 : _GEN_777; // @[Cat.scala 29:58]
  wire [7:0] _GEN_779 = 10'hff == pc[9:0] ? 8'h0 : _GEN_778; // @[Cat.scala 29:58]
  wire [7:0] _GEN_780 = 10'h100 == pc[9:0] ? 8'he3 : _GEN_779; // @[Cat.scala 29:58]
  wire [7:0] _GEN_781 = 10'h101 == pc[9:0] ? 8'h8c : _GEN_780; // @[Cat.scala 29:58]
  wire [7:0] _GEN_782 = 10'h102 == pc[9:0] ? 8'h7 : _GEN_781; // @[Cat.scala 29:58]
  wire [7:0] _GEN_783 = 10'h103 == pc[9:0] ? 8'hfe : _GEN_782; // @[Cat.scala 29:58]
  wire [7:0] _GEN_784 = 10'h104 == pc[9:0] ? 8'hef : _GEN_783; // @[Cat.scala 29:58]
  wire [7:0] _GEN_785 = 10'h105 == pc[9:0] ? 8'hf0 : _GEN_784; // @[Cat.scala 29:58]
  wire [7:0] _GEN_786 = 10'h106 == pc[9:0] ? 8'h5f : _GEN_785; // @[Cat.scala 29:58]
  wire [7:0] _GEN_787 = 10'h107 == pc[9:0] ? 8'hf1 : _GEN_786; // @[Cat.scala 29:58]
  wire [7:0] _GEN_788 = 10'h108 == pc[9:0] ? 8'h93 : _GEN_787; // @[Cat.scala 29:58]
  wire [7:0] _GEN_789 = 10'h109 == pc[9:0] ? 8'h7 : _GEN_788; // @[Cat.scala 29:58]
  wire [7:0] _GEN_790 = 10'h10a == pc[9:0] ? 8'h5 : _GEN_789; // @[Cat.scala 29:58]
  wire [7:0] _GEN_791 = 10'h10b == pc[9:0] ? 8'h0 : _GEN_790; // @[Cat.scala 29:58]
  wire [7:0] _GEN_792 = 10'h10c == pc[9:0] ? 8'h13 : _GEN_791; // @[Cat.scala 29:58]
  wire [7:0] _GEN_793 = 10'h10d == pc[9:0] ? 8'h85 : _GEN_792; // @[Cat.scala 29:58]
  wire [7:0] _GEN_794 = 10'h10e == pc[9:0] ? 8'h7 : _GEN_793; // @[Cat.scala 29:58]
  wire [7:0] _GEN_795 = 10'h10f == pc[9:0] ? 8'h0 : _GEN_794; // @[Cat.scala 29:58]
  wire [7:0] _GEN_796 = 10'h110 == pc[9:0] ? 8'hef : _GEN_795; // @[Cat.scala 29:58]
  wire [7:0] _GEN_797 = 10'h111 == pc[9:0] ? 8'hf0 : _GEN_796; // @[Cat.scala 29:58]
  wire [7:0] _GEN_798 = 10'h112 == pc[9:0] ? 8'h9f : _GEN_797; // @[Cat.scala 29:58]
  wire [7:0] _GEN_799 = 10'h113 == pc[9:0] ? 8'hf6 : _GEN_798; // @[Cat.scala 29:58]
  wire [7:0] _GEN_800 = 10'h114 == pc[9:0] ? 8'h23 : _GEN_799; // @[Cat.scala 29:58]
  wire [7:0] _GEN_801 = 10'h115 == pc[9:0] ? 8'h26 : _GEN_800; // @[Cat.scala 29:58]
  wire [7:0] _GEN_802 = 10'h116 == pc[9:0] ? 8'h4 : _GEN_801; // @[Cat.scala 29:58]
  wire [7:0] _GEN_803 = 10'h117 == pc[9:0] ? 8'hfe : _GEN_802; // @[Cat.scala 29:58]
  wire [7:0] _GEN_804 = 10'h118 == pc[9:0] ? 8'h6f : _GEN_803; // @[Cat.scala 29:58]
  wire [7:0] _GEN_805 = 10'h119 == pc[9:0] ? 8'h0 : _GEN_804; // @[Cat.scala 29:58]
  wire [7:0] _GEN_806 = 10'h11a == pc[9:0] ? 8'h0 : _GEN_805; // @[Cat.scala 29:58]
  wire [7:0] _GEN_807 = 10'h11b == pc[9:0] ? 8'h1 : _GEN_806; // @[Cat.scala 29:58]
  wire [7:0] _GEN_808 = 10'h11c == pc[9:0] ? 8'h83 : _GEN_807; // @[Cat.scala 29:58]
  wire [7:0] _GEN_809 = 10'h11d == pc[9:0] ? 8'h27 : _GEN_808; // @[Cat.scala 29:58]
  wire [7:0] _GEN_810 = 10'h11e == pc[9:0] ? 8'hc4 : _GEN_809; // @[Cat.scala 29:58]
  wire [7:0] _GEN_811 = 10'h11f == pc[9:0] ? 8'hfe : _GEN_810; // @[Cat.scala 29:58]
  wire [7:0] _GEN_812 = 10'h120 == pc[9:0] ? 8'h93 : _GEN_811; // @[Cat.scala 29:58]
  wire [7:0] _GEN_813 = 10'h121 == pc[9:0] ? 8'h87 : _GEN_812; // @[Cat.scala 29:58]
  wire [7:0] _GEN_814 = 10'h122 == pc[9:0] ? 8'h17 : _GEN_813; // @[Cat.scala 29:58]
  wire [7:0] _GEN_815 = 10'h123 == pc[9:0] ? 8'h0 : _GEN_814; // @[Cat.scala 29:58]
  wire [7:0] _GEN_816 = 10'h124 == pc[9:0] ? 8'h23 : _GEN_815; // @[Cat.scala 29:58]
  wire [7:0] _GEN_817 = 10'h125 == pc[9:0] ? 8'h26 : _GEN_816; // @[Cat.scala 29:58]
  wire [7:0] _GEN_818 = 10'h126 == pc[9:0] ? 8'hf4 : _GEN_817; // @[Cat.scala 29:58]
  wire [7:0] _GEN_819 = 10'h127 == pc[9:0] ? 8'hfe : _GEN_818; // @[Cat.scala 29:58]
  wire [7:0] _GEN_820 = 10'h128 == pc[9:0] ? 8'h3 : _GEN_819; // @[Cat.scala 29:58]
  wire [7:0] _GEN_821 = 10'h129 == pc[9:0] ? 8'h27 : _GEN_820; // @[Cat.scala 29:58]
  wire [7:0] _GEN_822 = 10'h12a == pc[9:0] ? 8'hc4 : _GEN_821; // @[Cat.scala 29:58]
  wire [7:0] _GEN_823 = 10'h12b == pc[9:0] ? 8'hfe : _GEN_822; // @[Cat.scala 29:58]
  wire [7:0] _GEN_824 = 10'h12c == pc[9:0] ? 8'hb7 : _GEN_823; // @[Cat.scala 29:58]
  wire [7:0] _GEN_825 = 10'h12d == pc[9:0] ? 8'h57 : _GEN_824; // @[Cat.scala 29:58]
  wire [7:0] _GEN_826 = 10'h12e == pc[9:0] ? 8'h89 : _GEN_825; // @[Cat.scala 29:58]
  wire [7:0] _GEN_827 = 10'h12f == pc[9:0] ? 8'h0 : _GEN_826; // @[Cat.scala 29:58]
  wire [7:0] _GEN_828 = 10'h130 == pc[9:0] ? 8'h93 : _GEN_827; // @[Cat.scala 29:58]
  wire [7:0] _GEN_829 = 10'h131 == pc[9:0] ? 8'h87 : _GEN_828; // @[Cat.scala 29:58]
  wire [7:0] _GEN_830 = 10'h132 == pc[9:0] ? 8'hf7 : _GEN_829; // @[Cat.scala 29:58]
  wire [7:0] _GEN_831 = 10'h133 == pc[9:0] ? 8'h43 : _GEN_830; // @[Cat.scala 29:58]
  wire [7:0] _GEN_832 = 10'h134 == pc[9:0] ? 8'he3 : _GEN_831; // @[Cat.scala 29:58]
  wire [7:0] _GEN_833 = 10'h135 == pc[9:0] ? 8'hd4 : _GEN_832; // @[Cat.scala 29:58]
  wire [7:0] _GEN_834 = 10'h136 == pc[9:0] ? 8'he7 : _GEN_833; // @[Cat.scala 29:58]
  wire [7:0] _GEN_835 = 10'h137 == pc[9:0] ? 8'hfe : _GEN_834; // @[Cat.scala 29:58]
  wire [7:0] _GEN_836 = 10'h138 == pc[9:0] ? 8'h13 : _GEN_835; // @[Cat.scala 29:58]
  wire [7:0] _GEN_837 = 10'h139 == pc[9:0] ? 8'h5 : _GEN_836; // @[Cat.scala 29:58]
  wire [7:0] _GEN_838 = 10'h13a == pc[9:0] ? 8'h0 : _GEN_837; // @[Cat.scala 29:58]
  wire [7:0] _GEN_839 = 10'h13b == pc[9:0] ? 8'h0 : _GEN_838; // @[Cat.scala 29:58]
  wire [7:0] _GEN_840 = 10'h13c == pc[9:0] ? 8'hef : _GEN_839; // @[Cat.scala 29:58]
  wire [7:0] _GEN_841 = 10'h13d == pc[9:0] ? 8'hf0 : _GEN_840; // @[Cat.scala 29:58]
  wire [7:0] _GEN_842 = 10'h13e == pc[9:0] ? 8'hdf : _GEN_841; // @[Cat.scala 29:58]
  wire [7:0] _GEN_843 = 10'h13f == pc[9:0] ? 8'hf3 : _GEN_842; // @[Cat.scala 29:58]
  wire [7:0] _GEN_844 = 10'h140 == pc[9:0] ? 8'h6f : _GEN_843; // @[Cat.scala 29:58]
  wire [7:0] _GEN_845 = 10'h141 == pc[9:0] ? 8'hf0 : _GEN_844; // @[Cat.scala 29:58]
  wire [7:0] _GEN_846 = 10'h142 == pc[9:0] ? 8'h9f : _GEN_845; // @[Cat.scala 29:58]
  wire [7:0] _GEN_847 = 10'h143 == pc[9:0] ? 8'hfb : _GEN_846; // @[Cat.scala 29:58]
  wire [7:0] _GEN_848 = 10'h144 == pc[9:0] ? 8'h0 : _GEN_847; // @[Cat.scala 29:58]
  wire [7:0] _GEN_849 = 10'h145 == pc[9:0] ? 8'h0 : _GEN_848; // @[Cat.scala 29:58]
  wire [7:0] _GEN_850 = 10'h146 == pc[9:0] ? 8'h0 : _GEN_849; // @[Cat.scala 29:58]
  wire [7:0] _GEN_851 = 10'h147 == pc[9:0] ? 8'h0 : _GEN_850; // @[Cat.scala 29:58]
  wire [7:0] _GEN_852 = 10'h148 == pc[9:0] ? 8'h0 : _GEN_851; // @[Cat.scala 29:58]
  wire [7:0] _GEN_853 = 10'h149 == pc[9:0] ? 8'h0 : _GEN_852; // @[Cat.scala 29:58]
  wire [7:0] _GEN_854 = 10'h14a == pc[9:0] ? 8'h0 : _GEN_853; // @[Cat.scala 29:58]
  wire [7:0] _GEN_855 = 10'h14b == pc[9:0] ? 8'h0 : _GEN_854; // @[Cat.scala 29:58]
  wire [7:0] _GEN_856 = 10'h14c == pc[9:0] ? 8'h0 : _GEN_855; // @[Cat.scala 29:58]
  wire [7:0] _GEN_857 = 10'h14d == pc[9:0] ? 8'h0 : _GEN_856; // @[Cat.scala 29:58]
  wire [7:0] _GEN_858 = 10'h14e == pc[9:0] ? 8'h0 : _GEN_857; // @[Cat.scala 29:58]
  wire [7:0] _GEN_859 = 10'h14f == pc[9:0] ? 8'h0 : _GEN_858; // @[Cat.scala 29:58]
  wire [7:0] _GEN_860 = 10'h150 == pc[9:0] ? 8'h0 : _GEN_859; // @[Cat.scala 29:58]
  wire [7:0] _GEN_861 = 10'h151 == pc[9:0] ? 8'h0 : _GEN_860; // @[Cat.scala 29:58]
  wire [7:0] _GEN_862 = 10'h152 == pc[9:0] ? 8'h0 : _GEN_861; // @[Cat.scala 29:58]
  wire [7:0] _GEN_863 = 10'h153 == pc[9:0] ? 8'h0 : _GEN_862; // @[Cat.scala 29:58]
  wire [7:0] _GEN_864 = 10'h154 == pc[9:0] ? 8'h0 : _GEN_863; // @[Cat.scala 29:58]
  wire [7:0] _GEN_865 = 10'h155 == pc[9:0] ? 8'h0 : _GEN_864; // @[Cat.scala 29:58]
  wire [7:0] _GEN_866 = 10'h156 == pc[9:0] ? 8'h0 : _GEN_865; // @[Cat.scala 29:58]
  wire [7:0] _GEN_867 = 10'h157 == pc[9:0] ? 8'h0 : _GEN_866; // @[Cat.scala 29:58]
  wire [7:0] _GEN_868 = 10'h158 == pc[9:0] ? 8'h0 : _GEN_867; // @[Cat.scala 29:58]
  wire [7:0] _GEN_869 = 10'h159 == pc[9:0] ? 8'h0 : _GEN_868; // @[Cat.scala 29:58]
  wire [7:0] _GEN_870 = 10'h15a == pc[9:0] ? 8'h0 : _GEN_869; // @[Cat.scala 29:58]
  wire [7:0] _GEN_871 = 10'h15b == pc[9:0] ? 8'h0 : _GEN_870; // @[Cat.scala 29:58]
  wire [7:0] _GEN_872 = 10'h15c == pc[9:0] ? 8'h0 : _GEN_871; // @[Cat.scala 29:58]
  wire [7:0] _GEN_873 = 10'h15d == pc[9:0] ? 8'h0 : _GEN_872; // @[Cat.scala 29:58]
  wire [7:0] _GEN_874 = 10'h15e == pc[9:0] ? 8'h0 : _GEN_873; // @[Cat.scala 29:58]
  wire [7:0] _GEN_875 = 10'h15f == pc[9:0] ? 8'h0 : _GEN_874; // @[Cat.scala 29:58]
  wire [7:0] _GEN_876 = 10'h160 == pc[9:0] ? 8'h0 : _GEN_875; // @[Cat.scala 29:58]
  wire [7:0] _GEN_877 = 10'h161 == pc[9:0] ? 8'h0 : _GEN_876; // @[Cat.scala 29:58]
  wire [7:0] _GEN_878 = 10'h162 == pc[9:0] ? 8'h0 : _GEN_877; // @[Cat.scala 29:58]
  wire [7:0] _GEN_879 = 10'h163 == pc[9:0] ? 8'h0 : _GEN_878; // @[Cat.scala 29:58]
  wire [7:0] _GEN_880 = 10'h164 == pc[9:0] ? 8'h0 : _GEN_879; // @[Cat.scala 29:58]
  wire [7:0] _GEN_881 = 10'h165 == pc[9:0] ? 8'h0 : _GEN_880; // @[Cat.scala 29:58]
  wire [7:0] _GEN_882 = 10'h166 == pc[9:0] ? 8'h0 : _GEN_881; // @[Cat.scala 29:58]
  wire [7:0] _GEN_883 = 10'h167 == pc[9:0] ? 8'h0 : _GEN_882; // @[Cat.scala 29:58]
  wire [7:0] _GEN_884 = 10'h168 == pc[9:0] ? 8'h0 : _GEN_883; // @[Cat.scala 29:58]
  wire [7:0] _GEN_885 = 10'h169 == pc[9:0] ? 8'h0 : _GEN_884; // @[Cat.scala 29:58]
  wire [7:0] _GEN_886 = 10'h16a == pc[9:0] ? 8'h0 : _GEN_885; // @[Cat.scala 29:58]
  wire [7:0] _GEN_887 = 10'h16b == pc[9:0] ? 8'h0 : _GEN_886; // @[Cat.scala 29:58]
  wire [7:0] _GEN_888 = 10'h16c == pc[9:0] ? 8'h0 : _GEN_887; // @[Cat.scala 29:58]
  wire [7:0] _GEN_889 = 10'h16d == pc[9:0] ? 8'h0 : _GEN_888; // @[Cat.scala 29:58]
  wire [7:0] _GEN_890 = 10'h16e == pc[9:0] ? 8'h0 : _GEN_889; // @[Cat.scala 29:58]
  wire [7:0] _GEN_891 = 10'h16f == pc[9:0] ? 8'h0 : _GEN_890; // @[Cat.scala 29:58]
  wire [7:0] _GEN_892 = 10'h170 == pc[9:0] ? 8'h0 : _GEN_891; // @[Cat.scala 29:58]
  wire [7:0] _GEN_893 = 10'h171 == pc[9:0] ? 8'h0 : _GEN_892; // @[Cat.scala 29:58]
  wire [7:0] _GEN_894 = 10'h172 == pc[9:0] ? 8'h0 : _GEN_893; // @[Cat.scala 29:58]
  wire [7:0] _GEN_895 = 10'h173 == pc[9:0] ? 8'h0 : _GEN_894; // @[Cat.scala 29:58]
  wire [7:0] _GEN_896 = 10'h174 == pc[9:0] ? 8'h0 : _GEN_895; // @[Cat.scala 29:58]
  wire [7:0] _GEN_897 = 10'h175 == pc[9:0] ? 8'h0 : _GEN_896; // @[Cat.scala 29:58]
  wire [7:0] _GEN_898 = 10'h176 == pc[9:0] ? 8'h0 : _GEN_897; // @[Cat.scala 29:58]
  wire [7:0] _GEN_899 = 10'h177 == pc[9:0] ? 8'h0 : _GEN_898; // @[Cat.scala 29:58]
  wire [7:0] _GEN_900 = 10'h178 == pc[9:0] ? 8'h0 : _GEN_899; // @[Cat.scala 29:58]
  wire [7:0] _GEN_901 = 10'h179 == pc[9:0] ? 8'h0 : _GEN_900; // @[Cat.scala 29:58]
  wire [7:0] _GEN_902 = 10'h17a == pc[9:0] ? 8'h0 : _GEN_901; // @[Cat.scala 29:58]
  wire [7:0] _GEN_903 = 10'h17b == pc[9:0] ? 8'h0 : _GEN_902; // @[Cat.scala 29:58]
  wire [7:0] _GEN_904 = 10'h17c == pc[9:0] ? 8'h0 : _GEN_903; // @[Cat.scala 29:58]
  wire [7:0] _GEN_905 = 10'h17d == pc[9:0] ? 8'h0 : _GEN_904; // @[Cat.scala 29:58]
  wire [7:0] _GEN_906 = 10'h17e == pc[9:0] ? 8'h0 : _GEN_905; // @[Cat.scala 29:58]
  wire [7:0] _GEN_907 = 10'h17f == pc[9:0] ? 8'h0 : _GEN_906; // @[Cat.scala 29:58]
  wire [7:0] _GEN_908 = 10'h180 == pc[9:0] ? 8'h0 : _GEN_907; // @[Cat.scala 29:58]
  wire [7:0] _GEN_909 = 10'h181 == pc[9:0] ? 8'h0 : _GEN_908; // @[Cat.scala 29:58]
  wire [7:0] _GEN_910 = 10'h182 == pc[9:0] ? 8'h0 : _GEN_909; // @[Cat.scala 29:58]
  wire [7:0] _GEN_911 = 10'h183 == pc[9:0] ? 8'h0 : _GEN_910; // @[Cat.scala 29:58]
  wire [7:0] _GEN_912 = 10'h184 == pc[9:0] ? 8'h0 : _GEN_911; // @[Cat.scala 29:58]
  wire [7:0] _GEN_913 = 10'h185 == pc[9:0] ? 8'h0 : _GEN_912; // @[Cat.scala 29:58]
  wire [7:0] _GEN_914 = 10'h186 == pc[9:0] ? 8'h0 : _GEN_913; // @[Cat.scala 29:58]
  wire [7:0] _GEN_915 = 10'h187 == pc[9:0] ? 8'h0 : _GEN_914; // @[Cat.scala 29:58]
  wire [7:0] _GEN_916 = 10'h188 == pc[9:0] ? 8'h0 : _GEN_915; // @[Cat.scala 29:58]
  wire [7:0] _GEN_917 = 10'h189 == pc[9:0] ? 8'h0 : _GEN_916; // @[Cat.scala 29:58]
  wire [7:0] _GEN_918 = 10'h18a == pc[9:0] ? 8'h0 : _GEN_917; // @[Cat.scala 29:58]
  wire [7:0] _GEN_919 = 10'h18b == pc[9:0] ? 8'h0 : _GEN_918; // @[Cat.scala 29:58]
  wire [7:0] _GEN_920 = 10'h18c == pc[9:0] ? 8'h0 : _GEN_919; // @[Cat.scala 29:58]
  wire [7:0] _GEN_921 = 10'h18d == pc[9:0] ? 8'h0 : _GEN_920; // @[Cat.scala 29:58]
  wire [7:0] _GEN_922 = 10'h18e == pc[9:0] ? 8'h0 : _GEN_921; // @[Cat.scala 29:58]
  wire [7:0] _GEN_923 = 10'h18f == pc[9:0] ? 8'h0 : _GEN_922; // @[Cat.scala 29:58]
  wire [7:0] _GEN_924 = 10'h190 == pc[9:0] ? 8'h0 : _GEN_923; // @[Cat.scala 29:58]
  wire [7:0] _GEN_925 = 10'h191 == pc[9:0] ? 8'h0 : _GEN_924; // @[Cat.scala 29:58]
  wire [7:0] _GEN_926 = 10'h192 == pc[9:0] ? 8'h0 : _GEN_925; // @[Cat.scala 29:58]
  wire [7:0] _GEN_927 = 10'h193 == pc[9:0] ? 8'h0 : _GEN_926; // @[Cat.scala 29:58]
  wire [7:0] _GEN_928 = 10'h194 == pc[9:0] ? 8'h0 : _GEN_927; // @[Cat.scala 29:58]
  wire [7:0] _GEN_929 = 10'h195 == pc[9:0] ? 8'h0 : _GEN_928; // @[Cat.scala 29:58]
  wire [7:0] _GEN_930 = 10'h196 == pc[9:0] ? 8'h0 : _GEN_929; // @[Cat.scala 29:58]
  wire [7:0] _GEN_931 = 10'h197 == pc[9:0] ? 8'h0 : _GEN_930; // @[Cat.scala 29:58]
  wire [7:0] _GEN_932 = 10'h198 == pc[9:0] ? 8'h0 : _GEN_931; // @[Cat.scala 29:58]
  wire [7:0] _GEN_933 = 10'h199 == pc[9:0] ? 8'h0 : _GEN_932; // @[Cat.scala 29:58]
  wire [7:0] _GEN_934 = 10'h19a == pc[9:0] ? 8'h0 : _GEN_933; // @[Cat.scala 29:58]
  wire [7:0] _GEN_935 = 10'h19b == pc[9:0] ? 8'h0 : _GEN_934; // @[Cat.scala 29:58]
  wire [7:0] _GEN_936 = 10'h19c == pc[9:0] ? 8'h0 : _GEN_935; // @[Cat.scala 29:58]
  wire [7:0] _GEN_937 = 10'h19d == pc[9:0] ? 8'h0 : _GEN_936; // @[Cat.scala 29:58]
  wire [7:0] _GEN_938 = 10'h19e == pc[9:0] ? 8'h0 : _GEN_937; // @[Cat.scala 29:58]
  wire [7:0] _GEN_939 = 10'h19f == pc[9:0] ? 8'h0 : _GEN_938; // @[Cat.scala 29:58]
  wire [7:0] _GEN_940 = 10'h1a0 == pc[9:0] ? 8'h0 : _GEN_939; // @[Cat.scala 29:58]
  wire [7:0] _GEN_941 = 10'h1a1 == pc[9:0] ? 8'h0 : _GEN_940; // @[Cat.scala 29:58]
  wire [7:0] _GEN_942 = 10'h1a2 == pc[9:0] ? 8'h0 : _GEN_941; // @[Cat.scala 29:58]
  wire [7:0] _GEN_943 = 10'h1a3 == pc[9:0] ? 8'h0 : _GEN_942; // @[Cat.scala 29:58]
  wire [7:0] _GEN_944 = 10'h1a4 == pc[9:0] ? 8'h0 : _GEN_943; // @[Cat.scala 29:58]
  wire [7:0] _GEN_945 = 10'h1a5 == pc[9:0] ? 8'h0 : _GEN_944; // @[Cat.scala 29:58]
  wire [7:0] _GEN_946 = 10'h1a6 == pc[9:0] ? 8'h0 : _GEN_945; // @[Cat.scala 29:58]
  wire [7:0] _GEN_947 = 10'h1a7 == pc[9:0] ? 8'h0 : _GEN_946; // @[Cat.scala 29:58]
  wire [7:0] _GEN_948 = 10'h1a8 == pc[9:0] ? 8'h0 : _GEN_947; // @[Cat.scala 29:58]
  wire [7:0] _GEN_949 = 10'h1a9 == pc[9:0] ? 8'h0 : _GEN_948; // @[Cat.scala 29:58]
  wire [7:0] _GEN_950 = 10'h1aa == pc[9:0] ? 8'h0 : _GEN_949; // @[Cat.scala 29:58]
  wire [7:0] _GEN_951 = 10'h1ab == pc[9:0] ? 8'h0 : _GEN_950; // @[Cat.scala 29:58]
  wire [7:0] _GEN_952 = 10'h1ac == pc[9:0] ? 8'h0 : _GEN_951; // @[Cat.scala 29:58]
  wire [7:0] _GEN_953 = 10'h1ad == pc[9:0] ? 8'h0 : _GEN_952; // @[Cat.scala 29:58]
  wire [7:0] _GEN_954 = 10'h1ae == pc[9:0] ? 8'h0 : _GEN_953; // @[Cat.scala 29:58]
  wire [7:0] _GEN_955 = 10'h1af == pc[9:0] ? 8'h0 : _GEN_954; // @[Cat.scala 29:58]
  wire [7:0] _GEN_956 = 10'h1b0 == pc[9:0] ? 8'h0 : _GEN_955; // @[Cat.scala 29:58]
  wire [7:0] _GEN_957 = 10'h1b1 == pc[9:0] ? 8'h0 : _GEN_956; // @[Cat.scala 29:58]
  wire [7:0] _GEN_958 = 10'h1b2 == pc[9:0] ? 8'h0 : _GEN_957; // @[Cat.scala 29:58]
  wire [7:0] _GEN_959 = 10'h1b3 == pc[9:0] ? 8'h0 : _GEN_958; // @[Cat.scala 29:58]
  wire [7:0] _GEN_960 = 10'h1b4 == pc[9:0] ? 8'h0 : _GEN_959; // @[Cat.scala 29:58]
  wire [7:0] _GEN_961 = 10'h1b5 == pc[9:0] ? 8'h0 : _GEN_960; // @[Cat.scala 29:58]
  wire [7:0] _GEN_962 = 10'h1b6 == pc[9:0] ? 8'h0 : _GEN_961; // @[Cat.scala 29:58]
  wire [7:0] _GEN_963 = 10'h1b7 == pc[9:0] ? 8'h0 : _GEN_962; // @[Cat.scala 29:58]
  wire [7:0] _GEN_964 = 10'h1b8 == pc[9:0] ? 8'h0 : _GEN_963; // @[Cat.scala 29:58]
  wire [7:0] _GEN_965 = 10'h1b9 == pc[9:0] ? 8'h0 : _GEN_964; // @[Cat.scala 29:58]
  wire [7:0] _GEN_966 = 10'h1ba == pc[9:0] ? 8'h0 : _GEN_965; // @[Cat.scala 29:58]
  wire [7:0] _GEN_967 = 10'h1bb == pc[9:0] ? 8'h0 : _GEN_966; // @[Cat.scala 29:58]
  wire [7:0] _GEN_968 = 10'h1bc == pc[9:0] ? 8'h0 : _GEN_967; // @[Cat.scala 29:58]
  wire [7:0] _GEN_969 = 10'h1bd == pc[9:0] ? 8'h0 : _GEN_968; // @[Cat.scala 29:58]
  wire [7:0] _GEN_970 = 10'h1be == pc[9:0] ? 8'h0 : _GEN_969; // @[Cat.scala 29:58]
  wire [7:0] _GEN_971 = 10'h1bf == pc[9:0] ? 8'h0 : _GEN_970; // @[Cat.scala 29:58]
  wire [7:0] _GEN_972 = 10'h1c0 == pc[9:0] ? 8'h0 : _GEN_971; // @[Cat.scala 29:58]
  wire [7:0] _GEN_973 = 10'h1c1 == pc[9:0] ? 8'h0 : _GEN_972; // @[Cat.scala 29:58]
  wire [7:0] _GEN_974 = 10'h1c2 == pc[9:0] ? 8'h0 : _GEN_973; // @[Cat.scala 29:58]
  wire [7:0] _GEN_975 = 10'h1c3 == pc[9:0] ? 8'h0 : _GEN_974; // @[Cat.scala 29:58]
  wire [7:0] _GEN_976 = 10'h1c4 == pc[9:0] ? 8'h0 : _GEN_975; // @[Cat.scala 29:58]
  wire [7:0] _GEN_977 = 10'h1c5 == pc[9:0] ? 8'h0 : _GEN_976; // @[Cat.scala 29:58]
  wire [7:0] _GEN_978 = 10'h1c6 == pc[9:0] ? 8'h0 : _GEN_977; // @[Cat.scala 29:58]
  wire [7:0] _GEN_979 = 10'h1c7 == pc[9:0] ? 8'h0 : _GEN_978; // @[Cat.scala 29:58]
  wire [7:0] _GEN_980 = 10'h1c8 == pc[9:0] ? 8'h0 : _GEN_979; // @[Cat.scala 29:58]
  wire [7:0] _GEN_981 = 10'h1c9 == pc[9:0] ? 8'h0 : _GEN_980; // @[Cat.scala 29:58]
  wire [7:0] _GEN_982 = 10'h1ca == pc[9:0] ? 8'h0 : _GEN_981; // @[Cat.scala 29:58]
  wire [7:0] _GEN_983 = 10'h1cb == pc[9:0] ? 8'h0 : _GEN_982; // @[Cat.scala 29:58]
  wire [7:0] _GEN_984 = 10'h1cc == pc[9:0] ? 8'h0 : _GEN_983; // @[Cat.scala 29:58]
  wire [7:0] _GEN_985 = 10'h1cd == pc[9:0] ? 8'h0 : _GEN_984; // @[Cat.scala 29:58]
  wire [7:0] _GEN_986 = 10'h1ce == pc[9:0] ? 8'h0 : _GEN_985; // @[Cat.scala 29:58]
  wire [7:0] _GEN_987 = 10'h1cf == pc[9:0] ? 8'h0 : _GEN_986; // @[Cat.scala 29:58]
  wire [7:0] _GEN_988 = 10'h1d0 == pc[9:0] ? 8'h0 : _GEN_987; // @[Cat.scala 29:58]
  wire [7:0] _GEN_989 = 10'h1d1 == pc[9:0] ? 8'h0 : _GEN_988; // @[Cat.scala 29:58]
  wire [7:0] _GEN_990 = 10'h1d2 == pc[9:0] ? 8'h0 : _GEN_989; // @[Cat.scala 29:58]
  wire [7:0] _GEN_991 = 10'h1d3 == pc[9:0] ? 8'h0 : _GEN_990; // @[Cat.scala 29:58]
  wire [7:0] _GEN_992 = 10'h1d4 == pc[9:0] ? 8'h0 : _GEN_991; // @[Cat.scala 29:58]
  wire [7:0] _GEN_993 = 10'h1d5 == pc[9:0] ? 8'h0 : _GEN_992; // @[Cat.scala 29:58]
  wire [7:0] _GEN_994 = 10'h1d6 == pc[9:0] ? 8'h0 : _GEN_993; // @[Cat.scala 29:58]
  wire [7:0] _GEN_995 = 10'h1d7 == pc[9:0] ? 8'h0 : _GEN_994; // @[Cat.scala 29:58]
  wire [7:0] _GEN_996 = 10'h1d8 == pc[9:0] ? 8'h0 : _GEN_995; // @[Cat.scala 29:58]
  wire [7:0] _GEN_997 = 10'h1d9 == pc[9:0] ? 8'h0 : _GEN_996; // @[Cat.scala 29:58]
  wire [7:0] _GEN_998 = 10'h1da == pc[9:0] ? 8'h0 : _GEN_997; // @[Cat.scala 29:58]
  wire [7:0] _GEN_999 = 10'h1db == pc[9:0] ? 8'h0 : _GEN_998; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1000 = 10'h1dc == pc[9:0] ? 8'h0 : _GEN_999; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1001 = 10'h1dd == pc[9:0] ? 8'h0 : _GEN_1000; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1002 = 10'h1de == pc[9:0] ? 8'h0 : _GEN_1001; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1003 = 10'h1df == pc[9:0] ? 8'h0 : _GEN_1002; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1004 = 10'h1e0 == pc[9:0] ? 8'h0 : _GEN_1003; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1005 = 10'h1e1 == pc[9:0] ? 8'h0 : _GEN_1004; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1006 = 10'h1e2 == pc[9:0] ? 8'h0 : _GEN_1005; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1007 = 10'h1e3 == pc[9:0] ? 8'h0 : _GEN_1006; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1008 = 10'h1e4 == pc[9:0] ? 8'h0 : _GEN_1007; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1009 = 10'h1e5 == pc[9:0] ? 8'h0 : _GEN_1008; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1010 = 10'h1e6 == pc[9:0] ? 8'h0 : _GEN_1009; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1011 = 10'h1e7 == pc[9:0] ? 8'h0 : _GEN_1010; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1012 = 10'h1e8 == pc[9:0] ? 8'h0 : _GEN_1011; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1013 = 10'h1e9 == pc[9:0] ? 8'h0 : _GEN_1012; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1014 = 10'h1ea == pc[9:0] ? 8'h0 : _GEN_1013; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1015 = 10'h1eb == pc[9:0] ? 8'h0 : _GEN_1014; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1016 = 10'h1ec == pc[9:0] ? 8'h0 : _GEN_1015; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1017 = 10'h1ed == pc[9:0] ? 8'h0 : _GEN_1016; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1018 = 10'h1ee == pc[9:0] ? 8'h0 : _GEN_1017; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1019 = 10'h1ef == pc[9:0] ? 8'h0 : _GEN_1018; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1020 = 10'h1f0 == pc[9:0] ? 8'h0 : _GEN_1019; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1021 = 10'h1f1 == pc[9:0] ? 8'h0 : _GEN_1020; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1022 = 10'h1f2 == pc[9:0] ? 8'h0 : _GEN_1021; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1023 = 10'h1f3 == pc[9:0] ? 8'h0 : _GEN_1022; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1024 = 10'h1f4 == pc[9:0] ? 8'h0 : _GEN_1023; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1025 = 10'h1f5 == pc[9:0] ? 8'h0 : _GEN_1024; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1026 = 10'h1f6 == pc[9:0] ? 8'h0 : _GEN_1025; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1027 = 10'h1f7 == pc[9:0] ? 8'h0 : _GEN_1026; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1028 = 10'h1f8 == pc[9:0] ? 8'h0 : _GEN_1027; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1029 = 10'h1f9 == pc[9:0] ? 8'h0 : _GEN_1028; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1030 = 10'h1fa == pc[9:0] ? 8'h0 : _GEN_1029; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1031 = 10'h1fb == pc[9:0] ? 8'h0 : _GEN_1030; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1032 = 10'h1fc == pc[9:0] ? 8'h0 : _GEN_1031; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1033 = 10'h1fd == pc[9:0] ? 8'h0 : _GEN_1032; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1034 = 10'h1fe == pc[9:0] ? 8'h0 : _GEN_1033; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1035 = 10'h1ff == pc[9:0] ? 8'h0 : _GEN_1034; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1036 = 10'h200 == pc[9:0] ? 8'h0 : _GEN_1035; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1037 = 10'h201 == pc[9:0] ? 8'h0 : _GEN_1036; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1038 = 10'h202 == pc[9:0] ? 8'h0 : _GEN_1037; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1039 = 10'h203 == pc[9:0] ? 8'h0 : _GEN_1038; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1040 = 10'h204 == pc[9:0] ? 8'h0 : _GEN_1039; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1041 = 10'h205 == pc[9:0] ? 8'h0 : _GEN_1040; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1042 = 10'h206 == pc[9:0] ? 8'h0 : _GEN_1041; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1043 = 10'h207 == pc[9:0] ? 8'h0 : _GEN_1042; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1044 = 10'h208 == pc[9:0] ? 8'h0 : _GEN_1043; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1045 = 10'h209 == pc[9:0] ? 8'h0 : _GEN_1044; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1046 = 10'h20a == pc[9:0] ? 8'h0 : _GEN_1045; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1047 = 10'h20b == pc[9:0] ? 8'h0 : _GEN_1046; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1049 = 10'h1 == _T_1[9:0] ? 8'h21 : 8'h97; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1050 = 10'h2 == _T_1[9:0] ? 8'h0 : _GEN_1049; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1051 = 10'h3 == _T_1[9:0] ? 8'h0 : _GEN_1050; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1052 = 10'h4 == _T_1[9:0] ? 8'h93 : _GEN_1051; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1053 = 10'h5 == _T_1[9:0] ? 8'h81 : _GEN_1052; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1054 = 10'h6 == _T_1[9:0] ? 8'h1 : _GEN_1053; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1055 = 10'h7 == _T_1[9:0] ? 8'h97 : _GEN_1054; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1056 = 10'h8 == _T_1[9:0] ? 8'h17 : _GEN_1055; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1057 = 10'h9 == _T_1[9:0] ? 8'h11 : _GEN_1056; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1058 = 10'ha == _T_1[9:0] ? 8'h0 : _GEN_1057; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1059 = 10'hb == _T_1[9:0] ? 8'h0 : _GEN_1058; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1060 = 10'hc == _T_1[9:0] ? 8'h13 : _GEN_1059; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1061 = 10'hd == _T_1[9:0] ? 8'h1 : _GEN_1060; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1062 = 10'he == _T_1[9:0] ? 8'h81 : _GEN_1061; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1063 = 10'hf == _T_1[9:0] ? 8'hff : _GEN_1062; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1064 = 10'h10 == _T_1[9:0] ? 8'h33 : _GEN_1063; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1065 = 10'h11 == _T_1[9:0] ? 8'h4 : _GEN_1064; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1066 = 10'h12 == _T_1[9:0] ? 8'h1 : _GEN_1065; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1067 = 10'h13 == _T_1[9:0] ? 8'h0 : _GEN_1066; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1068 = 10'h14 == _T_1[9:0] ? 8'h6f : _GEN_1067; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1069 = 10'h15 == _T_1[9:0] ? 8'h0 : _GEN_1068; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1070 = 10'h16 == _T_1[9:0] ? 8'h80 : _GEN_1069; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1071 = 10'h17 == _T_1[9:0] ? 8'h9 : _GEN_1070; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1072 = 10'h18 == _T_1[9:0] ? 8'h13 : _GEN_1071; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1073 = 10'h19 == _T_1[9:0] ? 8'h1 : _GEN_1072; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1074 = 10'h1a == _T_1[9:0] ? 8'h1 : _GEN_1073; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1075 = 10'h1b == _T_1[9:0] ? 8'hfe : _GEN_1074; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1076 = 10'h1c == _T_1[9:0] ? 8'h23 : _GEN_1075; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1077 = 10'h1d == _T_1[9:0] ? 8'h2e : _GEN_1076; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1078 = 10'h1e == _T_1[9:0] ? 8'h81 : _GEN_1077; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1079 = 10'h1f == _T_1[9:0] ? 8'h0 : _GEN_1078; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1080 = 10'h20 == _T_1[9:0] ? 8'h13 : _GEN_1079; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1081 = 10'h21 == _T_1[9:0] ? 8'h4 : _GEN_1080; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1082 = 10'h22 == _T_1[9:0] ? 8'h1 : _GEN_1081; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1083 = 10'h23 == _T_1[9:0] ? 8'h2 : _GEN_1082; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1084 = 10'h24 == _T_1[9:0] ? 8'hb7 : _GEN_1083; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1085 = 10'h25 == _T_1[9:0] ? 8'h27 : _GEN_1084; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1086 = 10'h26 == _T_1[9:0] ? 8'h0 : _GEN_1085; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1087 = 10'h27 == _T_1[9:0] ? 8'h0 : _GEN_1086; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1088 = 10'h28 == _T_1[9:0] ? 8'h93 : _GEN_1087; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1089 = 10'h29 == _T_1[9:0] ? 8'h87 : _GEN_1088; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1090 = 10'h2a == _T_1[9:0] ? 8'h7 : _GEN_1089; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1091 = 10'h2b == _T_1[9:0] ? 8'h20 : _GEN_1090; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1092 = 10'h2c == _T_1[9:0] ? 8'h23 : _GEN_1091; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1093 = 10'h2d == _T_1[9:0] ? 8'h26 : _GEN_1092; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1094 = 10'h2e == _T_1[9:0] ? 8'hf4 : _GEN_1093; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1095 = 10'h2f == _T_1[9:0] ? 8'hfe : _GEN_1094; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1096 = 10'h30 == _T_1[9:0] ? 8'h83 : _GEN_1095; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1097 = 10'h31 == _T_1[9:0] ? 8'h27 : _GEN_1096; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1098 = 10'h32 == _T_1[9:0] ? 8'hc4 : _GEN_1097; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1099 = 10'h33 == _T_1[9:0] ? 8'hfe : _GEN_1098; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1100 = 10'h34 == _T_1[9:0] ? 8'h83 : _GEN_1099; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1101 = 10'h35 == _T_1[9:0] ? 8'ha7 : _GEN_1100; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1102 = 10'h36 == _T_1[9:0] ? 8'h7 : _GEN_1101; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1103 = 10'h37 == _T_1[9:0] ? 8'h0 : _GEN_1102; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1104 = 10'h38 == _T_1[9:0] ? 8'h13 : _GEN_1103; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1105 = 10'h39 == _T_1[9:0] ? 8'h85 : _GEN_1104; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1106 = 10'h3a == _T_1[9:0] ? 8'h7 : _GEN_1105; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1107 = 10'h3b == _T_1[9:0] ? 8'h0 : _GEN_1106; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1108 = 10'h3c == _T_1[9:0] ? 8'h3 : _GEN_1107; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1109 = 10'h3d == _T_1[9:0] ? 8'h24 : _GEN_1108; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1110 = 10'h3e == _T_1[9:0] ? 8'hc1 : _GEN_1109; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1111 = 10'h3f == _T_1[9:0] ? 8'h1 : _GEN_1110; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1112 = 10'h40 == _T_1[9:0] ? 8'h13 : _GEN_1111; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1113 = 10'h41 == _T_1[9:0] ? 8'h1 : _GEN_1112; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1114 = 10'h42 == _T_1[9:0] ? 8'h1 : _GEN_1113; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1115 = 10'h43 == _T_1[9:0] ? 8'h2 : _GEN_1114; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1116 = 10'h44 == _T_1[9:0] ? 8'h67 : _GEN_1115; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1117 = 10'h45 == _T_1[9:0] ? 8'h80 : _GEN_1116; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1118 = 10'h46 == _T_1[9:0] ? 8'h0 : _GEN_1117; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1119 = 10'h47 == _T_1[9:0] ? 8'h0 : _GEN_1118; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1120 = 10'h48 == _T_1[9:0] ? 8'h13 : _GEN_1119; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1121 = 10'h49 == _T_1[9:0] ? 8'h1 : _GEN_1120; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1122 = 10'h4a == _T_1[9:0] ? 8'h1 : _GEN_1121; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1123 = 10'h4b == _T_1[9:0] ? 8'hfe : _GEN_1122; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1124 = 10'h4c == _T_1[9:0] ? 8'h23 : _GEN_1123; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1125 = 10'h4d == _T_1[9:0] ? 8'h2e : _GEN_1124; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1126 = 10'h4e == _T_1[9:0] ? 8'h81 : _GEN_1125; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1127 = 10'h4f == _T_1[9:0] ? 8'h0 : _GEN_1126; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1128 = 10'h50 == _T_1[9:0] ? 8'h13 : _GEN_1127; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1129 = 10'h51 == _T_1[9:0] ? 8'h4 : _GEN_1128; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1130 = 10'h52 == _T_1[9:0] ? 8'h1 : _GEN_1129; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1131 = 10'h53 == _T_1[9:0] ? 8'h2 : _GEN_1130; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1132 = 10'h54 == _T_1[9:0] ? 8'hb7 : _GEN_1131; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1133 = 10'h55 == _T_1[9:0] ? 8'h27 : _GEN_1132; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1134 = 10'h56 == _T_1[9:0] ? 8'h0 : _GEN_1133; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1135 = 10'h57 == _T_1[9:0] ? 8'h0 : _GEN_1134; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1136 = 10'h58 == _T_1[9:0] ? 8'h93 : _GEN_1135; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1137 = 10'h59 == _T_1[9:0] ? 8'h87 : _GEN_1136; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1138 = 10'h5a == _T_1[9:0] ? 8'h7 : _GEN_1137; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1139 = 10'h5b == _T_1[9:0] ? 8'h10 : _GEN_1138; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1140 = 10'h5c == _T_1[9:0] ? 8'h23 : _GEN_1139; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1141 = 10'h5d == _T_1[9:0] ? 8'h26 : _GEN_1140; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1142 = 10'h5e == _T_1[9:0] ? 8'hf4 : _GEN_1141; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1143 = 10'h5f == _T_1[9:0] ? 8'hfe : _GEN_1142; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1144 = 10'h60 == _T_1[9:0] ? 8'h83 : _GEN_1143; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1145 = 10'h61 == _T_1[9:0] ? 8'h27 : _GEN_1144; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1146 = 10'h62 == _T_1[9:0] ? 8'hc4 : _GEN_1145; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1147 = 10'h63 == _T_1[9:0] ? 8'hfe : _GEN_1146; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1148 = 10'h64 == _T_1[9:0] ? 8'h83 : _GEN_1147; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1149 = 10'h65 == _T_1[9:0] ? 8'ha7 : _GEN_1148; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1150 = 10'h66 == _T_1[9:0] ? 8'h7 : _GEN_1149; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1151 = 10'h67 == _T_1[9:0] ? 8'h0 : _GEN_1150; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1152 = 10'h68 == _T_1[9:0] ? 8'h13 : _GEN_1151; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1153 = 10'h69 == _T_1[9:0] ? 8'h85 : _GEN_1152; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1154 = 10'h6a == _T_1[9:0] ? 8'h7 : _GEN_1153; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1155 = 10'h6b == _T_1[9:0] ? 8'h0 : _GEN_1154; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1156 = 10'h6c == _T_1[9:0] ? 8'h3 : _GEN_1155; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1157 = 10'h6d == _T_1[9:0] ? 8'h24 : _GEN_1156; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1158 = 10'h6e == _T_1[9:0] ? 8'hc1 : _GEN_1157; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1159 = 10'h6f == _T_1[9:0] ? 8'h1 : _GEN_1158; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1160 = 10'h70 == _T_1[9:0] ? 8'h13 : _GEN_1159; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1161 = 10'h71 == _T_1[9:0] ? 8'h1 : _GEN_1160; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1162 = 10'h72 == _T_1[9:0] ? 8'h1 : _GEN_1161; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1163 = 10'h73 == _T_1[9:0] ? 8'h2 : _GEN_1162; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1164 = 10'h74 == _T_1[9:0] ? 8'h67 : _GEN_1163; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1165 = 10'h75 == _T_1[9:0] ? 8'h80 : _GEN_1164; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1166 = 10'h76 == _T_1[9:0] ? 8'h0 : _GEN_1165; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1167 = 10'h77 == _T_1[9:0] ? 8'h0 : _GEN_1166; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1168 = 10'h78 == _T_1[9:0] ? 8'h13 : _GEN_1167; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1169 = 10'h79 == _T_1[9:0] ? 8'h1 : _GEN_1168; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1170 = 10'h7a == _T_1[9:0] ? 8'h1 : _GEN_1169; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1171 = 10'h7b == _T_1[9:0] ? 8'hfd : _GEN_1170; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1172 = 10'h7c == _T_1[9:0] ? 8'h23 : _GEN_1171; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1173 = 10'h7d == _T_1[9:0] ? 8'h26 : _GEN_1172; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1174 = 10'h7e == _T_1[9:0] ? 8'h81 : _GEN_1173; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1175 = 10'h7f == _T_1[9:0] ? 8'h2 : _GEN_1174; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1176 = 10'h80 == _T_1[9:0] ? 8'h13 : _GEN_1175; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1177 = 10'h81 == _T_1[9:0] ? 8'h4 : _GEN_1176; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1178 = 10'h82 == _T_1[9:0] ? 8'h1 : _GEN_1177; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1179 = 10'h83 == _T_1[9:0] ? 8'h3 : _GEN_1178; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1180 = 10'h84 == _T_1[9:0] ? 8'h23 : _GEN_1179; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1181 = 10'h85 == _T_1[9:0] ? 8'h2e : _GEN_1180; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1182 = 10'h86 == _T_1[9:0] ? 8'ha4 : _GEN_1181; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1183 = 10'h87 == _T_1[9:0] ? 8'hfc : _GEN_1182; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1184 = 10'h88 == _T_1[9:0] ? 8'hb7 : _GEN_1183; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1185 = 10'h89 == _T_1[9:0] ? 8'h27 : _GEN_1184; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1186 = 10'h8a == _T_1[9:0] ? 8'h0 : _GEN_1185; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1187 = 10'h8b == _T_1[9:0] ? 8'h0 : _GEN_1186; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1188 = 10'h8c == _T_1[9:0] ? 8'h23 : _GEN_1187; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1189 = 10'h8d == _T_1[9:0] ? 8'h26 : _GEN_1188; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1190 = 10'h8e == _T_1[9:0] ? 8'hf4 : _GEN_1189; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1191 = 10'h8f == _T_1[9:0] ? 8'hfe : _GEN_1190; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1192 = 10'h90 == _T_1[9:0] ? 8'h83 : _GEN_1191; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1193 = 10'h91 == _T_1[9:0] ? 8'h27 : _GEN_1192; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1194 = 10'h92 == _T_1[9:0] ? 8'hc4 : _GEN_1193; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1195 = 10'h93 == _T_1[9:0] ? 8'hfe : _GEN_1194; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1196 = 10'h94 == _T_1[9:0] ? 8'h3 : _GEN_1195; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1197 = 10'h95 == _T_1[9:0] ? 8'h27 : _GEN_1196; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1198 = 10'h96 == _T_1[9:0] ? 8'hc4 : _GEN_1197; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1199 = 10'h97 == _T_1[9:0] ? 8'hfd : _GEN_1198; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1200 = 10'h98 == _T_1[9:0] ? 8'h23 : _GEN_1199; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1201 = 10'h99 == _T_1[9:0] ? 8'ha0 : _GEN_1200; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1202 = 10'h9a == _T_1[9:0] ? 8'he7 : _GEN_1201; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1203 = 10'h9b == _T_1[9:0] ? 8'h0 : _GEN_1202; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1204 = 10'h9c == _T_1[9:0] ? 8'h13 : _GEN_1203; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1205 = 10'h9d == _T_1[9:0] ? 8'h0 : _GEN_1204; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1206 = 10'h9e == _T_1[9:0] ? 8'h0 : _GEN_1205; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1207 = 10'h9f == _T_1[9:0] ? 8'h0 : _GEN_1206; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1208 = 10'ha0 == _T_1[9:0] ? 8'h3 : _GEN_1207; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1209 = 10'ha1 == _T_1[9:0] ? 8'h24 : _GEN_1208; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1210 = 10'ha2 == _T_1[9:0] ? 8'hc1 : _GEN_1209; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1211 = 10'ha3 == _T_1[9:0] ? 8'h2 : _GEN_1210; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1212 = 10'ha4 == _T_1[9:0] ? 8'h13 : _GEN_1211; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1213 = 10'ha5 == _T_1[9:0] ? 8'h1 : _GEN_1212; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1214 = 10'ha6 == _T_1[9:0] ? 8'h1 : _GEN_1213; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1215 = 10'ha7 == _T_1[9:0] ? 8'h3 : _GEN_1214; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1216 = 10'ha8 == _T_1[9:0] ? 8'h67 : _GEN_1215; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1217 = 10'ha9 == _T_1[9:0] ? 8'h80 : _GEN_1216; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1218 = 10'haa == _T_1[9:0] ? 8'h0 : _GEN_1217; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1219 = 10'hab == _T_1[9:0] ? 8'h0 : _GEN_1218; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1220 = 10'hac == _T_1[9:0] ? 8'h13 : _GEN_1219; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1221 = 10'had == _T_1[9:0] ? 8'h1 : _GEN_1220; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1222 = 10'hae == _T_1[9:0] ? 8'h1 : _GEN_1221; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1223 = 10'haf == _T_1[9:0] ? 8'hfe : _GEN_1222; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1224 = 10'hb0 == _T_1[9:0] ? 8'h23 : _GEN_1223; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1225 = 10'hb1 == _T_1[9:0] ? 8'h2e : _GEN_1224; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1226 = 10'hb2 == _T_1[9:0] ? 8'h11 : _GEN_1225; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1227 = 10'hb3 == _T_1[9:0] ? 8'h0 : _GEN_1226; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1228 = 10'hb4 == _T_1[9:0] ? 8'h23 : _GEN_1227; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1229 = 10'hb5 == _T_1[9:0] ? 8'h2c : _GEN_1228; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1230 = 10'hb6 == _T_1[9:0] ? 8'h81 : _GEN_1229; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1231 = 10'hb7 == _T_1[9:0] ? 8'h0 : _GEN_1230; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1232 = 10'hb8 == _T_1[9:0] ? 8'h13 : _GEN_1231; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1233 = 10'hb9 == _T_1[9:0] ? 8'h4 : _GEN_1232; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1234 = 10'hba == _T_1[9:0] ? 8'h1 : _GEN_1233; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1235 = 10'hbb == _T_1[9:0] ? 8'h2 : _GEN_1234; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1236 = 10'hbc == _T_1[9:0] ? 8'h23 : _GEN_1235; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1237 = 10'hbd == _T_1[9:0] ? 8'h26 : _GEN_1236; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1238 = 10'hbe == _T_1[9:0] ? 8'h4 : _GEN_1237; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1239 = 10'hbf == _T_1[9:0] ? 8'hfe : _GEN_1238; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1240 = 10'hc0 == _T_1[9:0] ? 8'hb7 : _GEN_1239; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1241 = 10'hc1 == _T_1[9:0] ? 8'hc7 : _GEN_1240; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1242 = 10'hc2 == _T_1[9:0] ? 8'h0 : _GEN_1241; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1243 = 10'hc3 == _T_1[9:0] ? 8'h0 : _GEN_1242; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1244 = 10'hc4 == _T_1[9:0] ? 8'h13 : _GEN_1243; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1245 = 10'hc5 == _T_1[9:0] ? 8'h85 : _GEN_1244; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1246 = 10'hc6 == _T_1[9:0] ? 8'hf7 : _GEN_1245; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1247 = 10'hc7 == _T_1[9:0] ? 8'hee : _GEN_1246; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1248 = 10'hc8 == _T_1[9:0] ? 8'hef : _GEN_1247; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1249 = 10'hc9 == _T_1[9:0] ? 8'hf0 : _GEN_1248; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1250 = 10'hca == _T_1[9:0] ? 8'h1f : _GEN_1249; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1251 = 10'hcb == _T_1[9:0] ? 8'hfb : _GEN_1250; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1252 = 10'hcc == _T_1[9:0] ? 8'h23 : _GEN_1251; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1253 = 10'hcd == _T_1[9:0] ? 8'h26 : _GEN_1252; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1254 = 10'hce == _T_1[9:0] ? 8'h4 : _GEN_1253; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1255 = 10'hcf == _T_1[9:0] ? 8'hfe : _GEN_1254; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1256 = 10'hd0 == _T_1[9:0] ? 8'h6f : _GEN_1255; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1257 = 10'hd1 == _T_1[9:0] ? 8'h0 : _GEN_1256; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1258 = 10'hd2 == _T_1[9:0] ? 8'h0 : _GEN_1257; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1259 = 10'hd3 == _T_1[9:0] ? 8'h1 : _GEN_1258; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1260 = 10'hd4 == _T_1[9:0] ? 8'h83 : _GEN_1259; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1261 = 10'hd5 == _T_1[9:0] ? 8'h27 : _GEN_1260; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1262 = 10'hd6 == _T_1[9:0] ? 8'hc4 : _GEN_1261; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1263 = 10'hd7 == _T_1[9:0] ? 8'hfe : _GEN_1262; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1264 = 10'hd8 == _T_1[9:0] ? 8'h93 : _GEN_1263; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1265 = 10'hd9 == _T_1[9:0] ? 8'h87 : _GEN_1264; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1266 = 10'hda == _T_1[9:0] ? 8'h17 : _GEN_1265; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1267 = 10'hdb == _T_1[9:0] ? 8'h0 : _GEN_1266; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1268 = 10'hdc == _T_1[9:0] ? 8'h23 : _GEN_1267; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1269 = 10'hdd == _T_1[9:0] ? 8'h26 : _GEN_1268; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1270 = 10'hde == _T_1[9:0] ? 8'hf4 : _GEN_1269; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1271 = 10'hdf == _T_1[9:0] ? 8'hfe : _GEN_1270; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1272 = 10'he0 == _T_1[9:0] ? 8'h3 : _GEN_1271; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1273 = 10'he1 == _T_1[9:0] ? 8'h27 : _GEN_1272; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1274 = 10'he2 == _T_1[9:0] ? 8'hc4 : _GEN_1273; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1275 = 10'he3 == _T_1[9:0] ? 8'hfe : _GEN_1274; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1276 = 10'he4 == _T_1[9:0] ? 8'hb7 : _GEN_1275; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1277 = 10'he5 == _T_1[9:0] ? 8'h17 : _GEN_1276; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1278 = 10'he6 == _T_1[9:0] ? 8'h7a : _GEN_1277; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1279 = 10'he7 == _T_1[9:0] ? 8'h0 : _GEN_1278; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1280 = 10'he8 == _T_1[9:0] ? 8'h93 : _GEN_1279; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1281 = 10'he9 == _T_1[9:0] ? 8'h87 : _GEN_1280; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1282 = 10'hea == _T_1[9:0] ? 8'hf7 : _GEN_1281; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1283 = 10'heb == _T_1[9:0] ? 8'h1f : _GEN_1282; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1284 = 10'hec == _T_1[9:0] ? 8'he3 : _GEN_1283; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1285 = 10'hed == _T_1[9:0] ? 8'hd4 : _GEN_1284; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1286 = 10'hee == _T_1[9:0] ? 8'he7 : _GEN_1285; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1287 = 10'hef == _T_1[9:0] ? 8'hfe : _GEN_1286; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1288 = 10'hf0 == _T_1[9:0] ? 8'h13 : _GEN_1287; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1289 = 10'hf1 == _T_1[9:0] ? 8'h5 : _GEN_1288; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1290 = 10'hf2 == _T_1[9:0] ? 8'h0 : _GEN_1289; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1291 = 10'hf3 == _T_1[9:0] ? 8'h0 : _GEN_1290; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1292 = 10'hf4 == _T_1[9:0] ? 8'hef : _GEN_1291; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1293 = 10'hf5 == _T_1[9:0] ? 8'hf0 : _GEN_1292; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1294 = 10'hf6 == _T_1[9:0] ? 8'h5f : _GEN_1293; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1295 = 10'hf7 == _T_1[9:0] ? 8'hf8 : _GEN_1294; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1296 = 10'hf8 == _T_1[9:0] ? 8'hef : _GEN_1295; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1297 = 10'hf9 == _T_1[9:0] ? 8'hf0 : _GEN_1296; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1298 = 10'hfa == _T_1[9:0] ? 8'h1f : _GEN_1297; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1299 = 10'hfb == _T_1[9:0] ? 8'hf5 : _GEN_1298; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1300 = 10'hfc == _T_1[9:0] ? 8'h93 : _GEN_1299; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1301 = 10'hfd == _T_1[9:0] ? 8'h7 : _GEN_1300; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1302 = 10'hfe == _T_1[9:0] ? 8'h5 : _GEN_1301; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1303 = 10'hff == _T_1[9:0] ? 8'h0 : _GEN_1302; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1304 = 10'h100 == _T_1[9:0] ? 8'he3 : _GEN_1303; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1305 = 10'h101 == _T_1[9:0] ? 8'h8c : _GEN_1304; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1306 = 10'h102 == _T_1[9:0] ? 8'h7 : _GEN_1305; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1307 = 10'h103 == _T_1[9:0] ? 8'hfe : _GEN_1306; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1308 = 10'h104 == _T_1[9:0] ? 8'hef : _GEN_1307; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1309 = 10'h105 == _T_1[9:0] ? 8'hf0 : _GEN_1308; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1310 = 10'h106 == _T_1[9:0] ? 8'h5f : _GEN_1309; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1311 = 10'h107 == _T_1[9:0] ? 8'hf1 : _GEN_1310; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1312 = 10'h108 == _T_1[9:0] ? 8'h93 : _GEN_1311; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1313 = 10'h109 == _T_1[9:0] ? 8'h7 : _GEN_1312; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1314 = 10'h10a == _T_1[9:0] ? 8'h5 : _GEN_1313; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1315 = 10'h10b == _T_1[9:0] ? 8'h0 : _GEN_1314; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1316 = 10'h10c == _T_1[9:0] ? 8'h13 : _GEN_1315; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1317 = 10'h10d == _T_1[9:0] ? 8'h85 : _GEN_1316; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1318 = 10'h10e == _T_1[9:0] ? 8'h7 : _GEN_1317; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1319 = 10'h10f == _T_1[9:0] ? 8'h0 : _GEN_1318; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1320 = 10'h110 == _T_1[9:0] ? 8'hef : _GEN_1319; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1321 = 10'h111 == _T_1[9:0] ? 8'hf0 : _GEN_1320; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1322 = 10'h112 == _T_1[9:0] ? 8'h9f : _GEN_1321; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1323 = 10'h113 == _T_1[9:0] ? 8'hf6 : _GEN_1322; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1324 = 10'h114 == _T_1[9:0] ? 8'h23 : _GEN_1323; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1325 = 10'h115 == _T_1[9:0] ? 8'h26 : _GEN_1324; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1326 = 10'h116 == _T_1[9:0] ? 8'h4 : _GEN_1325; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1327 = 10'h117 == _T_1[9:0] ? 8'hfe : _GEN_1326; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1328 = 10'h118 == _T_1[9:0] ? 8'h6f : _GEN_1327; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1329 = 10'h119 == _T_1[9:0] ? 8'h0 : _GEN_1328; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1330 = 10'h11a == _T_1[9:0] ? 8'h0 : _GEN_1329; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1331 = 10'h11b == _T_1[9:0] ? 8'h1 : _GEN_1330; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1332 = 10'h11c == _T_1[9:0] ? 8'h83 : _GEN_1331; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1333 = 10'h11d == _T_1[9:0] ? 8'h27 : _GEN_1332; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1334 = 10'h11e == _T_1[9:0] ? 8'hc4 : _GEN_1333; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1335 = 10'h11f == _T_1[9:0] ? 8'hfe : _GEN_1334; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1336 = 10'h120 == _T_1[9:0] ? 8'h93 : _GEN_1335; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1337 = 10'h121 == _T_1[9:0] ? 8'h87 : _GEN_1336; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1338 = 10'h122 == _T_1[9:0] ? 8'h17 : _GEN_1337; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1339 = 10'h123 == _T_1[9:0] ? 8'h0 : _GEN_1338; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1340 = 10'h124 == _T_1[9:0] ? 8'h23 : _GEN_1339; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1341 = 10'h125 == _T_1[9:0] ? 8'h26 : _GEN_1340; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1342 = 10'h126 == _T_1[9:0] ? 8'hf4 : _GEN_1341; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1343 = 10'h127 == _T_1[9:0] ? 8'hfe : _GEN_1342; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1344 = 10'h128 == _T_1[9:0] ? 8'h3 : _GEN_1343; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1345 = 10'h129 == _T_1[9:0] ? 8'h27 : _GEN_1344; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1346 = 10'h12a == _T_1[9:0] ? 8'hc4 : _GEN_1345; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1347 = 10'h12b == _T_1[9:0] ? 8'hfe : _GEN_1346; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1348 = 10'h12c == _T_1[9:0] ? 8'hb7 : _GEN_1347; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1349 = 10'h12d == _T_1[9:0] ? 8'h57 : _GEN_1348; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1350 = 10'h12e == _T_1[9:0] ? 8'h89 : _GEN_1349; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1351 = 10'h12f == _T_1[9:0] ? 8'h0 : _GEN_1350; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1352 = 10'h130 == _T_1[9:0] ? 8'h93 : _GEN_1351; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1353 = 10'h131 == _T_1[9:0] ? 8'h87 : _GEN_1352; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1354 = 10'h132 == _T_1[9:0] ? 8'hf7 : _GEN_1353; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1355 = 10'h133 == _T_1[9:0] ? 8'h43 : _GEN_1354; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1356 = 10'h134 == _T_1[9:0] ? 8'he3 : _GEN_1355; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1357 = 10'h135 == _T_1[9:0] ? 8'hd4 : _GEN_1356; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1358 = 10'h136 == _T_1[9:0] ? 8'he7 : _GEN_1357; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1359 = 10'h137 == _T_1[9:0] ? 8'hfe : _GEN_1358; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1360 = 10'h138 == _T_1[9:0] ? 8'h13 : _GEN_1359; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1361 = 10'h139 == _T_1[9:0] ? 8'h5 : _GEN_1360; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1362 = 10'h13a == _T_1[9:0] ? 8'h0 : _GEN_1361; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1363 = 10'h13b == _T_1[9:0] ? 8'h0 : _GEN_1362; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1364 = 10'h13c == _T_1[9:0] ? 8'hef : _GEN_1363; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1365 = 10'h13d == _T_1[9:0] ? 8'hf0 : _GEN_1364; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1366 = 10'h13e == _T_1[9:0] ? 8'hdf : _GEN_1365; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1367 = 10'h13f == _T_1[9:0] ? 8'hf3 : _GEN_1366; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1368 = 10'h140 == _T_1[9:0] ? 8'h6f : _GEN_1367; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1369 = 10'h141 == _T_1[9:0] ? 8'hf0 : _GEN_1368; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1370 = 10'h142 == _T_1[9:0] ? 8'h9f : _GEN_1369; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1371 = 10'h143 == _T_1[9:0] ? 8'hfb : _GEN_1370; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1372 = 10'h144 == _T_1[9:0] ? 8'h0 : _GEN_1371; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1373 = 10'h145 == _T_1[9:0] ? 8'h0 : _GEN_1372; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1374 = 10'h146 == _T_1[9:0] ? 8'h0 : _GEN_1373; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1375 = 10'h147 == _T_1[9:0] ? 8'h0 : _GEN_1374; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1376 = 10'h148 == _T_1[9:0] ? 8'h0 : _GEN_1375; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1377 = 10'h149 == _T_1[9:0] ? 8'h0 : _GEN_1376; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1378 = 10'h14a == _T_1[9:0] ? 8'h0 : _GEN_1377; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1379 = 10'h14b == _T_1[9:0] ? 8'h0 : _GEN_1378; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1380 = 10'h14c == _T_1[9:0] ? 8'h0 : _GEN_1379; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1381 = 10'h14d == _T_1[9:0] ? 8'h0 : _GEN_1380; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1382 = 10'h14e == _T_1[9:0] ? 8'h0 : _GEN_1381; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1383 = 10'h14f == _T_1[9:0] ? 8'h0 : _GEN_1382; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1384 = 10'h150 == _T_1[9:0] ? 8'h0 : _GEN_1383; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1385 = 10'h151 == _T_1[9:0] ? 8'h0 : _GEN_1384; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1386 = 10'h152 == _T_1[9:0] ? 8'h0 : _GEN_1385; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1387 = 10'h153 == _T_1[9:0] ? 8'h0 : _GEN_1386; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1388 = 10'h154 == _T_1[9:0] ? 8'h0 : _GEN_1387; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1389 = 10'h155 == _T_1[9:0] ? 8'h0 : _GEN_1388; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1390 = 10'h156 == _T_1[9:0] ? 8'h0 : _GEN_1389; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1391 = 10'h157 == _T_1[9:0] ? 8'h0 : _GEN_1390; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1392 = 10'h158 == _T_1[9:0] ? 8'h0 : _GEN_1391; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1393 = 10'h159 == _T_1[9:0] ? 8'h0 : _GEN_1392; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1394 = 10'h15a == _T_1[9:0] ? 8'h0 : _GEN_1393; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1395 = 10'h15b == _T_1[9:0] ? 8'h0 : _GEN_1394; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1396 = 10'h15c == _T_1[9:0] ? 8'h0 : _GEN_1395; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1397 = 10'h15d == _T_1[9:0] ? 8'h0 : _GEN_1396; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1398 = 10'h15e == _T_1[9:0] ? 8'h0 : _GEN_1397; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1399 = 10'h15f == _T_1[9:0] ? 8'h0 : _GEN_1398; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1400 = 10'h160 == _T_1[9:0] ? 8'h0 : _GEN_1399; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1401 = 10'h161 == _T_1[9:0] ? 8'h0 : _GEN_1400; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1402 = 10'h162 == _T_1[9:0] ? 8'h0 : _GEN_1401; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1403 = 10'h163 == _T_1[9:0] ? 8'h0 : _GEN_1402; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1404 = 10'h164 == _T_1[9:0] ? 8'h0 : _GEN_1403; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1405 = 10'h165 == _T_1[9:0] ? 8'h0 : _GEN_1404; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1406 = 10'h166 == _T_1[9:0] ? 8'h0 : _GEN_1405; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1407 = 10'h167 == _T_1[9:0] ? 8'h0 : _GEN_1406; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1408 = 10'h168 == _T_1[9:0] ? 8'h0 : _GEN_1407; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1409 = 10'h169 == _T_1[9:0] ? 8'h0 : _GEN_1408; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1410 = 10'h16a == _T_1[9:0] ? 8'h0 : _GEN_1409; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1411 = 10'h16b == _T_1[9:0] ? 8'h0 : _GEN_1410; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1412 = 10'h16c == _T_1[9:0] ? 8'h0 : _GEN_1411; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1413 = 10'h16d == _T_1[9:0] ? 8'h0 : _GEN_1412; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1414 = 10'h16e == _T_1[9:0] ? 8'h0 : _GEN_1413; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1415 = 10'h16f == _T_1[9:0] ? 8'h0 : _GEN_1414; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1416 = 10'h170 == _T_1[9:0] ? 8'h0 : _GEN_1415; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1417 = 10'h171 == _T_1[9:0] ? 8'h0 : _GEN_1416; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1418 = 10'h172 == _T_1[9:0] ? 8'h0 : _GEN_1417; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1419 = 10'h173 == _T_1[9:0] ? 8'h0 : _GEN_1418; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1420 = 10'h174 == _T_1[9:0] ? 8'h0 : _GEN_1419; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1421 = 10'h175 == _T_1[9:0] ? 8'h0 : _GEN_1420; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1422 = 10'h176 == _T_1[9:0] ? 8'h0 : _GEN_1421; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1423 = 10'h177 == _T_1[9:0] ? 8'h0 : _GEN_1422; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1424 = 10'h178 == _T_1[9:0] ? 8'h0 : _GEN_1423; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1425 = 10'h179 == _T_1[9:0] ? 8'h0 : _GEN_1424; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1426 = 10'h17a == _T_1[9:0] ? 8'h0 : _GEN_1425; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1427 = 10'h17b == _T_1[9:0] ? 8'h0 : _GEN_1426; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1428 = 10'h17c == _T_1[9:0] ? 8'h0 : _GEN_1427; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1429 = 10'h17d == _T_1[9:0] ? 8'h0 : _GEN_1428; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1430 = 10'h17e == _T_1[9:0] ? 8'h0 : _GEN_1429; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1431 = 10'h17f == _T_1[9:0] ? 8'h0 : _GEN_1430; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1432 = 10'h180 == _T_1[9:0] ? 8'h0 : _GEN_1431; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1433 = 10'h181 == _T_1[9:0] ? 8'h0 : _GEN_1432; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1434 = 10'h182 == _T_1[9:0] ? 8'h0 : _GEN_1433; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1435 = 10'h183 == _T_1[9:0] ? 8'h0 : _GEN_1434; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1436 = 10'h184 == _T_1[9:0] ? 8'h0 : _GEN_1435; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1437 = 10'h185 == _T_1[9:0] ? 8'h0 : _GEN_1436; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1438 = 10'h186 == _T_1[9:0] ? 8'h0 : _GEN_1437; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1439 = 10'h187 == _T_1[9:0] ? 8'h0 : _GEN_1438; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1440 = 10'h188 == _T_1[9:0] ? 8'h0 : _GEN_1439; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1441 = 10'h189 == _T_1[9:0] ? 8'h0 : _GEN_1440; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1442 = 10'h18a == _T_1[9:0] ? 8'h0 : _GEN_1441; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1443 = 10'h18b == _T_1[9:0] ? 8'h0 : _GEN_1442; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1444 = 10'h18c == _T_1[9:0] ? 8'h0 : _GEN_1443; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1445 = 10'h18d == _T_1[9:0] ? 8'h0 : _GEN_1444; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1446 = 10'h18e == _T_1[9:0] ? 8'h0 : _GEN_1445; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1447 = 10'h18f == _T_1[9:0] ? 8'h0 : _GEN_1446; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1448 = 10'h190 == _T_1[9:0] ? 8'h0 : _GEN_1447; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1449 = 10'h191 == _T_1[9:0] ? 8'h0 : _GEN_1448; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1450 = 10'h192 == _T_1[9:0] ? 8'h0 : _GEN_1449; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1451 = 10'h193 == _T_1[9:0] ? 8'h0 : _GEN_1450; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1452 = 10'h194 == _T_1[9:0] ? 8'h0 : _GEN_1451; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1453 = 10'h195 == _T_1[9:0] ? 8'h0 : _GEN_1452; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1454 = 10'h196 == _T_1[9:0] ? 8'h0 : _GEN_1453; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1455 = 10'h197 == _T_1[9:0] ? 8'h0 : _GEN_1454; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1456 = 10'h198 == _T_1[9:0] ? 8'h0 : _GEN_1455; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1457 = 10'h199 == _T_1[9:0] ? 8'h0 : _GEN_1456; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1458 = 10'h19a == _T_1[9:0] ? 8'h0 : _GEN_1457; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1459 = 10'h19b == _T_1[9:0] ? 8'h0 : _GEN_1458; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1460 = 10'h19c == _T_1[9:0] ? 8'h0 : _GEN_1459; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1461 = 10'h19d == _T_1[9:0] ? 8'h0 : _GEN_1460; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1462 = 10'h19e == _T_1[9:0] ? 8'h0 : _GEN_1461; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1463 = 10'h19f == _T_1[9:0] ? 8'h0 : _GEN_1462; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1464 = 10'h1a0 == _T_1[9:0] ? 8'h0 : _GEN_1463; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1465 = 10'h1a1 == _T_1[9:0] ? 8'h0 : _GEN_1464; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1466 = 10'h1a2 == _T_1[9:0] ? 8'h0 : _GEN_1465; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1467 = 10'h1a3 == _T_1[9:0] ? 8'h0 : _GEN_1466; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1468 = 10'h1a4 == _T_1[9:0] ? 8'h0 : _GEN_1467; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1469 = 10'h1a5 == _T_1[9:0] ? 8'h0 : _GEN_1468; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1470 = 10'h1a6 == _T_1[9:0] ? 8'h0 : _GEN_1469; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1471 = 10'h1a7 == _T_1[9:0] ? 8'h0 : _GEN_1470; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1472 = 10'h1a8 == _T_1[9:0] ? 8'h0 : _GEN_1471; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1473 = 10'h1a9 == _T_1[9:0] ? 8'h0 : _GEN_1472; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1474 = 10'h1aa == _T_1[9:0] ? 8'h0 : _GEN_1473; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1475 = 10'h1ab == _T_1[9:0] ? 8'h0 : _GEN_1474; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1476 = 10'h1ac == _T_1[9:0] ? 8'h0 : _GEN_1475; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1477 = 10'h1ad == _T_1[9:0] ? 8'h0 : _GEN_1476; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1478 = 10'h1ae == _T_1[9:0] ? 8'h0 : _GEN_1477; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1479 = 10'h1af == _T_1[9:0] ? 8'h0 : _GEN_1478; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1480 = 10'h1b0 == _T_1[9:0] ? 8'h0 : _GEN_1479; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1481 = 10'h1b1 == _T_1[9:0] ? 8'h0 : _GEN_1480; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1482 = 10'h1b2 == _T_1[9:0] ? 8'h0 : _GEN_1481; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1483 = 10'h1b3 == _T_1[9:0] ? 8'h0 : _GEN_1482; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1484 = 10'h1b4 == _T_1[9:0] ? 8'h0 : _GEN_1483; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1485 = 10'h1b5 == _T_1[9:0] ? 8'h0 : _GEN_1484; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1486 = 10'h1b6 == _T_1[9:0] ? 8'h0 : _GEN_1485; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1487 = 10'h1b7 == _T_1[9:0] ? 8'h0 : _GEN_1486; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1488 = 10'h1b8 == _T_1[9:0] ? 8'h0 : _GEN_1487; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1489 = 10'h1b9 == _T_1[9:0] ? 8'h0 : _GEN_1488; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1490 = 10'h1ba == _T_1[9:0] ? 8'h0 : _GEN_1489; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1491 = 10'h1bb == _T_1[9:0] ? 8'h0 : _GEN_1490; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1492 = 10'h1bc == _T_1[9:0] ? 8'h0 : _GEN_1491; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1493 = 10'h1bd == _T_1[9:0] ? 8'h0 : _GEN_1492; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1494 = 10'h1be == _T_1[9:0] ? 8'h0 : _GEN_1493; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1495 = 10'h1bf == _T_1[9:0] ? 8'h0 : _GEN_1494; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1496 = 10'h1c0 == _T_1[9:0] ? 8'h0 : _GEN_1495; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1497 = 10'h1c1 == _T_1[9:0] ? 8'h0 : _GEN_1496; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1498 = 10'h1c2 == _T_1[9:0] ? 8'h0 : _GEN_1497; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1499 = 10'h1c3 == _T_1[9:0] ? 8'h0 : _GEN_1498; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1500 = 10'h1c4 == _T_1[9:0] ? 8'h0 : _GEN_1499; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1501 = 10'h1c5 == _T_1[9:0] ? 8'h0 : _GEN_1500; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1502 = 10'h1c6 == _T_1[9:0] ? 8'h0 : _GEN_1501; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1503 = 10'h1c7 == _T_1[9:0] ? 8'h0 : _GEN_1502; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1504 = 10'h1c8 == _T_1[9:0] ? 8'h0 : _GEN_1503; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1505 = 10'h1c9 == _T_1[9:0] ? 8'h0 : _GEN_1504; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1506 = 10'h1ca == _T_1[9:0] ? 8'h0 : _GEN_1505; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1507 = 10'h1cb == _T_1[9:0] ? 8'h0 : _GEN_1506; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1508 = 10'h1cc == _T_1[9:0] ? 8'h0 : _GEN_1507; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1509 = 10'h1cd == _T_1[9:0] ? 8'h0 : _GEN_1508; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1510 = 10'h1ce == _T_1[9:0] ? 8'h0 : _GEN_1509; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1511 = 10'h1cf == _T_1[9:0] ? 8'h0 : _GEN_1510; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1512 = 10'h1d0 == _T_1[9:0] ? 8'h0 : _GEN_1511; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1513 = 10'h1d1 == _T_1[9:0] ? 8'h0 : _GEN_1512; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1514 = 10'h1d2 == _T_1[9:0] ? 8'h0 : _GEN_1513; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1515 = 10'h1d3 == _T_1[9:0] ? 8'h0 : _GEN_1514; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1516 = 10'h1d4 == _T_1[9:0] ? 8'h0 : _GEN_1515; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1517 = 10'h1d5 == _T_1[9:0] ? 8'h0 : _GEN_1516; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1518 = 10'h1d6 == _T_1[9:0] ? 8'h0 : _GEN_1517; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1519 = 10'h1d7 == _T_1[9:0] ? 8'h0 : _GEN_1518; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1520 = 10'h1d8 == _T_1[9:0] ? 8'h0 : _GEN_1519; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1521 = 10'h1d9 == _T_1[9:0] ? 8'h0 : _GEN_1520; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1522 = 10'h1da == _T_1[9:0] ? 8'h0 : _GEN_1521; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1523 = 10'h1db == _T_1[9:0] ? 8'h0 : _GEN_1522; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1524 = 10'h1dc == _T_1[9:0] ? 8'h0 : _GEN_1523; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1525 = 10'h1dd == _T_1[9:0] ? 8'h0 : _GEN_1524; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1526 = 10'h1de == _T_1[9:0] ? 8'h0 : _GEN_1525; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1527 = 10'h1df == _T_1[9:0] ? 8'h0 : _GEN_1526; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1528 = 10'h1e0 == _T_1[9:0] ? 8'h0 : _GEN_1527; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1529 = 10'h1e1 == _T_1[9:0] ? 8'h0 : _GEN_1528; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1530 = 10'h1e2 == _T_1[9:0] ? 8'h0 : _GEN_1529; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1531 = 10'h1e3 == _T_1[9:0] ? 8'h0 : _GEN_1530; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1532 = 10'h1e4 == _T_1[9:0] ? 8'h0 : _GEN_1531; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1533 = 10'h1e5 == _T_1[9:0] ? 8'h0 : _GEN_1532; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1534 = 10'h1e6 == _T_1[9:0] ? 8'h0 : _GEN_1533; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1535 = 10'h1e7 == _T_1[9:0] ? 8'h0 : _GEN_1534; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1536 = 10'h1e8 == _T_1[9:0] ? 8'h0 : _GEN_1535; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1537 = 10'h1e9 == _T_1[9:0] ? 8'h0 : _GEN_1536; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1538 = 10'h1ea == _T_1[9:0] ? 8'h0 : _GEN_1537; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1539 = 10'h1eb == _T_1[9:0] ? 8'h0 : _GEN_1538; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1540 = 10'h1ec == _T_1[9:0] ? 8'h0 : _GEN_1539; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1541 = 10'h1ed == _T_1[9:0] ? 8'h0 : _GEN_1540; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1542 = 10'h1ee == _T_1[9:0] ? 8'h0 : _GEN_1541; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1543 = 10'h1ef == _T_1[9:0] ? 8'h0 : _GEN_1542; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1544 = 10'h1f0 == _T_1[9:0] ? 8'h0 : _GEN_1543; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1545 = 10'h1f1 == _T_1[9:0] ? 8'h0 : _GEN_1544; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1546 = 10'h1f2 == _T_1[9:0] ? 8'h0 : _GEN_1545; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1547 = 10'h1f3 == _T_1[9:0] ? 8'h0 : _GEN_1546; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1548 = 10'h1f4 == _T_1[9:0] ? 8'h0 : _GEN_1547; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1549 = 10'h1f5 == _T_1[9:0] ? 8'h0 : _GEN_1548; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1550 = 10'h1f6 == _T_1[9:0] ? 8'h0 : _GEN_1549; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1551 = 10'h1f7 == _T_1[9:0] ? 8'h0 : _GEN_1550; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1552 = 10'h1f8 == _T_1[9:0] ? 8'h0 : _GEN_1551; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1553 = 10'h1f9 == _T_1[9:0] ? 8'h0 : _GEN_1552; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1554 = 10'h1fa == _T_1[9:0] ? 8'h0 : _GEN_1553; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1555 = 10'h1fb == _T_1[9:0] ? 8'h0 : _GEN_1554; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1556 = 10'h1fc == _T_1[9:0] ? 8'h0 : _GEN_1555; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1557 = 10'h1fd == _T_1[9:0] ? 8'h0 : _GEN_1556; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1558 = 10'h1fe == _T_1[9:0] ? 8'h0 : _GEN_1557; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1559 = 10'h1ff == _T_1[9:0] ? 8'h0 : _GEN_1558; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1560 = 10'h200 == _T_1[9:0] ? 8'h0 : _GEN_1559; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1561 = 10'h201 == _T_1[9:0] ? 8'h0 : _GEN_1560; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1562 = 10'h202 == _T_1[9:0] ? 8'h0 : _GEN_1561; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1563 = 10'h203 == _T_1[9:0] ? 8'h0 : _GEN_1562; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1564 = 10'h204 == _T_1[9:0] ? 8'h0 : _GEN_1563; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1565 = 10'h205 == _T_1[9:0] ? 8'h0 : _GEN_1564; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1566 = 10'h206 == _T_1[9:0] ? 8'h0 : _GEN_1565; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1567 = 10'h207 == _T_1[9:0] ? 8'h0 : _GEN_1566; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1568 = 10'h208 == _T_1[9:0] ? 8'h0 : _GEN_1567; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1569 = 10'h209 == _T_1[9:0] ? 8'h0 : _GEN_1568; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1570 = 10'h20a == _T_1[9:0] ? 8'h0 : _GEN_1569; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1571 = 10'h20b == _T_1[9:0] ? 8'h0 : _GEN_1570; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1573 = 10'h1 == _T_4[9:0] ? 8'h21 : 8'h97; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1574 = 10'h2 == _T_4[9:0] ? 8'h0 : _GEN_1573; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1575 = 10'h3 == _T_4[9:0] ? 8'h0 : _GEN_1574; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1576 = 10'h4 == _T_4[9:0] ? 8'h93 : _GEN_1575; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1577 = 10'h5 == _T_4[9:0] ? 8'h81 : _GEN_1576; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1578 = 10'h6 == _T_4[9:0] ? 8'h1 : _GEN_1577; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1579 = 10'h7 == _T_4[9:0] ? 8'h97 : _GEN_1578; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1580 = 10'h8 == _T_4[9:0] ? 8'h17 : _GEN_1579; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1581 = 10'h9 == _T_4[9:0] ? 8'h11 : _GEN_1580; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1582 = 10'ha == _T_4[9:0] ? 8'h0 : _GEN_1581; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1583 = 10'hb == _T_4[9:0] ? 8'h0 : _GEN_1582; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1584 = 10'hc == _T_4[9:0] ? 8'h13 : _GEN_1583; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1585 = 10'hd == _T_4[9:0] ? 8'h1 : _GEN_1584; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1586 = 10'he == _T_4[9:0] ? 8'h81 : _GEN_1585; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1587 = 10'hf == _T_4[9:0] ? 8'hff : _GEN_1586; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1588 = 10'h10 == _T_4[9:0] ? 8'h33 : _GEN_1587; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1589 = 10'h11 == _T_4[9:0] ? 8'h4 : _GEN_1588; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1590 = 10'h12 == _T_4[9:0] ? 8'h1 : _GEN_1589; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1591 = 10'h13 == _T_4[9:0] ? 8'h0 : _GEN_1590; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1592 = 10'h14 == _T_4[9:0] ? 8'h6f : _GEN_1591; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1593 = 10'h15 == _T_4[9:0] ? 8'h0 : _GEN_1592; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1594 = 10'h16 == _T_4[9:0] ? 8'h80 : _GEN_1593; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1595 = 10'h17 == _T_4[9:0] ? 8'h9 : _GEN_1594; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1596 = 10'h18 == _T_4[9:0] ? 8'h13 : _GEN_1595; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1597 = 10'h19 == _T_4[9:0] ? 8'h1 : _GEN_1596; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1598 = 10'h1a == _T_4[9:0] ? 8'h1 : _GEN_1597; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1599 = 10'h1b == _T_4[9:0] ? 8'hfe : _GEN_1598; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1600 = 10'h1c == _T_4[9:0] ? 8'h23 : _GEN_1599; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1601 = 10'h1d == _T_4[9:0] ? 8'h2e : _GEN_1600; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1602 = 10'h1e == _T_4[9:0] ? 8'h81 : _GEN_1601; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1603 = 10'h1f == _T_4[9:0] ? 8'h0 : _GEN_1602; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1604 = 10'h20 == _T_4[9:0] ? 8'h13 : _GEN_1603; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1605 = 10'h21 == _T_4[9:0] ? 8'h4 : _GEN_1604; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1606 = 10'h22 == _T_4[9:0] ? 8'h1 : _GEN_1605; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1607 = 10'h23 == _T_4[9:0] ? 8'h2 : _GEN_1606; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1608 = 10'h24 == _T_4[9:0] ? 8'hb7 : _GEN_1607; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1609 = 10'h25 == _T_4[9:0] ? 8'h27 : _GEN_1608; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1610 = 10'h26 == _T_4[9:0] ? 8'h0 : _GEN_1609; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1611 = 10'h27 == _T_4[9:0] ? 8'h0 : _GEN_1610; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1612 = 10'h28 == _T_4[9:0] ? 8'h93 : _GEN_1611; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1613 = 10'h29 == _T_4[9:0] ? 8'h87 : _GEN_1612; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1614 = 10'h2a == _T_4[9:0] ? 8'h7 : _GEN_1613; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1615 = 10'h2b == _T_4[9:0] ? 8'h20 : _GEN_1614; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1616 = 10'h2c == _T_4[9:0] ? 8'h23 : _GEN_1615; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1617 = 10'h2d == _T_4[9:0] ? 8'h26 : _GEN_1616; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1618 = 10'h2e == _T_4[9:0] ? 8'hf4 : _GEN_1617; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1619 = 10'h2f == _T_4[9:0] ? 8'hfe : _GEN_1618; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1620 = 10'h30 == _T_4[9:0] ? 8'h83 : _GEN_1619; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1621 = 10'h31 == _T_4[9:0] ? 8'h27 : _GEN_1620; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1622 = 10'h32 == _T_4[9:0] ? 8'hc4 : _GEN_1621; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1623 = 10'h33 == _T_4[9:0] ? 8'hfe : _GEN_1622; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1624 = 10'h34 == _T_4[9:0] ? 8'h83 : _GEN_1623; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1625 = 10'h35 == _T_4[9:0] ? 8'ha7 : _GEN_1624; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1626 = 10'h36 == _T_4[9:0] ? 8'h7 : _GEN_1625; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1627 = 10'h37 == _T_4[9:0] ? 8'h0 : _GEN_1626; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1628 = 10'h38 == _T_4[9:0] ? 8'h13 : _GEN_1627; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1629 = 10'h39 == _T_4[9:0] ? 8'h85 : _GEN_1628; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1630 = 10'h3a == _T_4[9:0] ? 8'h7 : _GEN_1629; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1631 = 10'h3b == _T_4[9:0] ? 8'h0 : _GEN_1630; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1632 = 10'h3c == _T_4[9:0] ? 8'h3 : _GEN_1631; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1633 = 10'h3d == _T_4[9:0] ? 8'h24 : _GEN_1632; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1634 = 10'h3e == _T_4[9:0] ? 8'hc1 : _GEN_1633; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1635 = 10'h3f == _T_4[9:0] ? 8'h1 : _GEN_1634; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1636 = 10'h40 == _T_4[9:0] ? 8'h13 : _GEN_1635; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1637 = 10'h41 == _T_4[9:0] ? 8'h1 : _GEN_1636; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1638 = 10'h42 == _T_4[9:0] ? 8'h1 : _GEN_1637; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1639 = 10'h43 == _T_4[9:0] ? 8'h2 : _GEN_1638; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1640 = 10'h44 == _T_4[9:0] ? 8'h67 : _GEN_1639; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1641 = 10'h45 == _T_4[9:0] ? 8'h80 : _GEN_1640; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1642 = 10'h46 == _T_4[9:0] ? 8'h0 : _GEN_1641; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1643 = 10'h47 == _T_4[9:0] ? 8'h0 : _GEN_1642; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1644 = 10'h48 == _T_4[9:0] ? 8'h13 : _GEN_1643; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1645 = 10'h49 == _T_4[9:0] ? 8'h1 : _GEN_1644; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1646 = 10'h4a == _T_4[9:0] ? 8'h1 : _GEN_1645; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1647 = 10'h4b == _T_4[9:0] ? 8'hfe : _GEN_1646; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1648 = 10'h4c == _T_4[9:0] ? 8'h23 : _GEN_1647; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1649 = 10'h4d == _T_4[9:0] ? 8'h2e : _GEN_1648; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1650 = 10'h4e == _T_4[9:0] ? 8'h81 : _GEN_1649; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1651 = 10'h4f == _T_4[9:0] ? 8'h0 : _GEN_1650; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1652 = 10'h50 == _T_4[9:0] ? 8'h13 : _GEN_1651; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1653 = 10'h51 == _T_4[9:0] ? 8'h4 : _GEN_1652; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1654 = 10'h52 == _T_4[9:0] ? 8'h1 : _GEN_1653; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1655 = 10'h53 == _T_4[9:0] ? 8'h2 : _GEN_1654; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1656 = 10'h54 == _T_4[9:0] ? 8'hb7 : _GEN_1655; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1657 = 10'h55 == _T_4[9:0] ? 8'h27 : _GEN_1656; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1658 = 10'h56 == _T_4[9:0] ? 8'h0 : _GEN_1657; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1659 = 10'h57 == _T_4[9:0] ? 8'h0 : _GEN_1658; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1660 = 10'h58 == _T_4[9:0] ? 8'h93 : _GEN_1659; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1661 = 10'h59 == _T_4[9:0] ? 8'h87 : _GEN_1660; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1662 = 10'h5a == _T_4[9:0] ? 8'h7 : _GEN_1661; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1663 = 10'h5b == _T_4[9:0] ? 8'h10 : _GEN_1662; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1664 = 10'h5c == _T_4[9:0] ? 8'h23 : _GEN_1663; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1665 = 10'h5d == _T_4[9:0] ? 8'h26 : _GEN_1664; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1666 = 10'h5e == _T_4[9:0] ? 8'hf4 : _GEN_1665; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1667 = 10'h5f == _T_4[9:0] ? 8'hfe : _GEN_1666; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1668 = 10'h60 == _T_4[9:0] ? 8'h83 : _GEN_1667; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1669 = 10'h61 == _T_4[9:0] ? 8'h27 : _GEN_1668; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1670 = 10'h62 == _T_4[9:0] ? 8'hc4 : _GEN_1669; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1671 = 10'h63 == _T_4[9:0] ? 8'hfe : _GEN_1670; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1672 = 10'h64 == _T_4[9:0] ? 8'h83 : _GEN_1671; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1673 = 10'h65 == _T_4[9:0] ? 8'ha7 : _GEN_1672; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1674 = 10'h66 == _T_4[9:0] ? 8'h7 : _GEN_1673; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1675 = 10'h67 == _T_4[9:0] ? 8'h0 : _GEN_1674; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1676 = 10'h68 == _T_4[9:0] ? 8'h13 : _GEN_1675; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1677 = 10'h69 == _T_4[9:0] ? 8'h85 : _GEN_1676; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1678 = 10'h6a == _T_4[9:0] ? 8'h7 : _GEN_1677; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1679 = 10'h6b == _T_4[9:0] ? 8'h0 : _GEN_1678; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1680 = 10'h6c == _T_4[9:0] ? 8'h3 : _GEN_1679; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1681 = 10'h6d == _T_4[9:0] ? 8'h24 : _GEN_1680; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1682 = 10'h6e == _T_4[9:0] ? 8'hc1 : _GEN_1681; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1683 = 10'h6f == _T_4[9:0] ? 8'h1 : _GEN_1682; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1684 = 10'h70 == _T_4[9:0] ? 8'h13 : _GEN_1683; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1685 = 10'h71 == _T_4[9:0] ? 8'h1 : _GEN_1684; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1686 = 10'h72 == _T_4[9:0] ? 8'h1 : _GEN_1685; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1687 = 10'h73 == _T_4[9:0] ? 8'h2 : _GEN_1686; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1688 = 10'h74 == _T_4[9:0] ? 8'h67 : _GEN_1687; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1689 = 10'h75 == _T_4[9:0] ? 8'h80 : _GEN_1688; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1690 = 10'h76 == _T_4[9:0] ? 8'h0 : _GEN_1689; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1691 = 10'h77 == _T_4[9:0] ? 8'h0 : _GEN_1690; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1692 = 10'h78 == _T_4[9:0] ? 8'h13 : _GEN_1691; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1693 = 10'h79 == _T_4[9:0] ? 8'h1 : _GEN_1692; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1694 = 10'h7a == _T_4[9:0] ? 8'h1 : _GEN_1693; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1695 = 10'h7b == _T_4[9:0] ? 8'hfd : _GEN_1694; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1696 = 10'h7c == _T_4[9:0] ? 8'h23 : _GEN_1695; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1697 = 10'h7d == _T_4[9:0] ? 8'h26 : _GEN_1696; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1698 = 10'h7e == _T_4[9:0] ? 8'h81 : _GEN_1697; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1699 = 10'h7f == _T_4[9:0] ? 8'h2 : _GEN_1698; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1700 = 10'h80 == _T_4[9:0] ? 8'h13 : _GEN_1699; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1701 = 10'h81 == _T_4[9:0] ? 8'h4 : _GEN_1700; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1702 = 10'h82 == _T_4[9:0] ? 8'h1 : _GEN_1701; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1703 = 10'h83 == _T_4[9:0] ? 8'h3 : _GEN_1702; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1704 = 10'h84 == _T_4[9:0] ? 8'h23 : _GEN_1703; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1705 = 10'h85 == _T_4[9:0] ? 8'h2e : _GEN_1704; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1706 = 10'h86 == _T_4[9:0] ? 8'ha4 : _GEN_1705; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1707 = 10'h87 == _T_4[9:0] ? 8'hfc : _GEN_1706; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1708 = 10'h88 == _T_4[9:0] ? 8'hb7 : _GEN_1707; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1709 = 10'h89 == _T_4[9:0] ? 8'h27 : _GEN_1708; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1710 = 10'h8a == _T_4[9:0] ? 8'h0 : _GEN_1709; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1711 = 10'h8b == _T_4[9:0] ? 8'h0 : _GEN_1710; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1712 = 10'h8c == _T_4[9:0] ? 8'h23 : _GEN_1711; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1713 = 10'h8d == _T_4[9:0] ? 8'h26 : _GEN_1712; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1714 = 10'h8e == _T_4[9:0] ? 8'hf4 : _GEN_1713; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1715 = 10'h8f == _T_4[9:0] ? 8'hfe : _GEN_1714; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1716 = 10'h90 == _T_4[9:0] ? 8'h83 : _GEN_1715; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1717 = 10'h91 == _T_4[9:0] ? 8'h27 : _GEN_1716; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1718 = 10'h92 == _T_4[9:0] ? 8'hc4 : _GEN_1717; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1719 = 10'h93 == _T_4[9:0] ? 8'hfe : _GEN_1718; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1720 = 10'h94 == _T_4[9:0] ? 8'h3 : _GEN_1719; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1721 = 10'h95 == _T_4[9:0] ? 8'h27 : _GEN_1720; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1722 = 10'h96 == _T_4[9:0] ? 8'hc4 : _GEN_1721; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1723 = 10'h97 == _T_4[9:0] ? 8'hfd : _GEN_1722; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1724 = 10'h98 == _T_4[9:0] ? 8'h23 : _GEN_1723; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1725 = 10'h99 == _T_4[9:0] ? 8'ha0 : _GEN_1724; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1726 = 10'h9a == _T_4[9:0] ? 8'he7 : _GEN_1725; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1727 = 10'h9b == _T_4[9:0] ? 8'h0 : _GEN_1726; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1728 = 10'h9c == _T_4[9:0] ? 8'h13 : _GEN_1727; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1729 = 10'h9d == _T_4[9:0] ? 8'h0 : _GEN_1728; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1730 = 10'h9e == _T_4[9:0] ? 8'h0 : _GEN_1729; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1731 = 10'h9f == _T_4[9:0] ? 8'h0 : _GEN_1730; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1732 = 10'ha0 == _T_4[9:0] ? 8'h3 : _GEN_1731; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1733 = 10'ha1 == _T_4[9:0] ? 8'h24 : _GEN_1732; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1734 = 10'ha2 == _T_4[9:0] ? 8'hc1 : _GEN_1733; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1735 = 10'ha3 == _T_4[9:0] ? 8'h2 : _GEN_1734; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1736 = 10'ha4 == _T_4[9:0] ? 8'h13 : _GEN_1735; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1737 = 10'ha5 == _T_4[9:0] ? 8'h1 : _GEN_1736; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1738 = 10'ha6 == _T_4[9:0] ? 8'h1 : _GEN_1737; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1739 = 10'ha7 == _T_4[9:0] ? 8'h3 : _GEN_1738; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1740 = 10'ha8 == _T_4[9:0] ? 8'h67 : _GEN_1739; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1741 = 10'ha9 == _T_4[9:0] ? 8'h80 : _GEN_1740; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1742 = 10'haa == _T_4[9:0] ? 8'h0 : _GEN_1741; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1743 = 10'hab == _T_4[9:0] ? 8'h0 : _GEN_1742; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1744 = 10'hac == _T_4[9:0] ? 8'h13 : _GEN_1743; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1745 = 10'had == _T_4[9:0] ? 8'h1 : _GEN_1744; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1746 = 10'hae == _T_4[9:0] ? 8'h1 : _GEN_1745; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1747 = 10'haf == _T_4[9:0] ? 8'hfe : _GEN_1746; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1748 = 10'hb0 == _T_4[9:0] ? 8'h23 : _GEN_1747; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1749 = 10'hb1 == _T_4[9:0] ? 8'h2e : _GEN_1748; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1750 = 10'hb2 == _T_4[9:0] ? 8'h11 : _GEN_1749; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1751 = 10'hb3 == _T_4[9:0] ? 8'h0 : _GEN_1750; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1752 = 10'hb4 == _T_4[9:0] ? 8'h23 : _GEN_1751; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1753 = 10'hb5 == _T_4[9:0] ? 8'h2c : _GEN_1752; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1754 = 10'hb6 == _T_4[9:0] ? 8'h81 : _GEN_1753; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1755 = 10'hb7 == _T_4[9:0] ? 8'h0 : _GEN_1754; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1756 = 10'hb8 == _T_4[9:0] ? 8'h13 : _GEN_1755; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1757 = 10'hb9 == _T_4[9:0] ? 8'h4 : _GEN_1756; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1758 = 10'hba == _T_4[9:0] ? 8'h1 : _GEN_1757; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1759 = 10'hbb == _T_4[9:0] ? 8'h2 : _GEN_1758; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1760 = 10'hbc == _T_4[9:0] ? 8'h23 : _GEN_1759; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1761 = 10'hbd == _T_4[9:0] ? 8'h26 : _GEN_1760; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1762 = 10'hbe == _T_4[9:0] ? 8'h4 : _GEN_1761; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1763 = 10'hbf == _T_4[9:0] ? 8'hfe : _GEN_1762; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1764 = 10'hc0 == _T_4[9:0] ? 8'hb7 : _GEN_1763; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1765 = 10'hc1 == _T_4[9:0] ? 8'hc7 : _GEN_1764; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1766 = 10'hc2 == _T_4[9:0] ? 8'h0 : _GEN_1765; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1767 = 10'hc3 == _T_4[9:0] ? 8'h0 : _GEN_1766; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1768 = 10'hc4 == _T_4[9:0] ? 8'h13 : _GEN_1767; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1769 = 10'hc5 == _T_4[9:0] ? 8'h85 : _GEN_1768; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1770 = 10'hc6 == _T_4[9:0] ? 8'hf7 : _GEN_1769; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1771 = 10'hc7 == _T_4[9:0] ? 8'hee : _GEN_1770; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1772 = 10'hc8 == _T_4[9:0] ? 8'hef : _GEN_1771; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1773 = 10'hc9 == _T_4[9:0] ? 8'hf0 : _GEN_1772; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1774 = 10'hca == _T_4[9:0] ? 8'h1f : _GEN_1773; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1775 = 10'hcb == _T_4[9:0] ? 8'hfb : _GEN_1774; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1776 = 10'hcc == _T_4[9:0] ? 8'h23 : _GEN_1775; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1777 = 10'hcd == _T_4[9:0] ? 8'h26 : _GEN_1776; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1778 = 10'hce == _T_4[9:0] ? 8'h4 : _GEN_1777; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1779 = 10'hcf == _T_4[9:0] ? 8'hfe : _GEN_1778; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1780 = 10'hd0 == _T_4[9:0] ? 8'h6f : _GEN_1779; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1781 = 10'hd1 == _T_4[9:0] ? 8'h0 : _GEN_1780; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1782 = 10'hd2 == _T_4[9:0] ? 8'h0 : _GEN_1781; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1783 = 10'hd3 == _T_4[9:0] ? 8'h1 : _GEN_1782; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1784 = 10'hd4 == _T_4[9:0] ? 8'h83 : _GEN_1783; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1785 = 10'hd5 == _T_4[9:0] ? 8'h27 : _GEN_1784; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1786 = 10'hd6 == _T_4[9:0] ? 8'hc4 : _GEN_1785; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1787 = 10'hd7 == _T_4[9:0] ? 8'hfe : _GEN_1786; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1788 = 10'hd8 == _T_4[9:0] ? 8'h93 : _GEN_1787; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1789 = 10'hd9 == _T_4[9:0] ? 8'h87 : _GEN_1788; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1790 = 10'hda == _T_4[9:0] ? 8'h17 : _GEN_1789; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1791 = 10'hdb == _T_4[9:0] ? 8'h0 : _GEN_1790; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1792 = 10'hdc == _T_4[9:0] ? 8'h23 : _GEN_1791; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1793 = 10'hdd == _T_4[9:0] ? 8'h26 : _GEN_1792; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1794 = 10'hde == _T_4[9:0] ? 8'hf4 : _GEN_1793; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1795 = 10'hdf == _T_4[9:0] ? 8'hfe : _GEN_1794; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1796 = 10'he0 == _T_4[9:0] ? 8'h3 : _GEN_1795; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1797 = 10'he1 == _T_4[9:0] ? 8'h27 : _GEN_1796; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1798 = 10'he2 == _T_4[9:0] ? 8'hc4 : _GEN_1797; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1799 = 10'he3 == _T_4[9:0] ? 8'hfe : _GEN_1798; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1800 = 10'he4 == _T_4[9:0] ? 8'hb7 : _GEN_1799; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1801 = 10'he5 == _T_4[9:0] ? 8'h17 : _GEN_1800; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1802 = 10'he6 == _T_4[9:0] ? 8'h7a : _GEN_1801; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1803 = 10'he7 == _T_4[9:0] ? 8'h0 : _GEN_1802; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1804 = 10'he8 == _T_4[9:0] ? 8'h93 : _GEN_1803; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1805 = 10'he9 == _T_4[9:0] ? 8'h87 : _GEN_1804; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1806 = 10'hea == _T_4[9:0] ? 8'hf7 : _GEN_1805; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1807 = 10'heb == _T_4[9:0] ? 8'h1f : _GEN_1806; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1808 = 10'hec == _T_4[9:0] ? 8'he3 : _GEN_1807; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1809 = 10'hed == _T_4[9:0] ? 8'hd4 : _GEN_1808; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1810 = 10'hee == _T_4[9:0] ? 8'he7 : _GEN_1809; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1811 = 10'hef == _T_4[9:0] ? 8'hfe : _GEN_1810; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1812 = 10'hf0 == _T_4[9:0] ? 8'h13 : _GEN_1811; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1813 = 10'hf1 == _T_4[9:0] ? 8'h5 : _GEN_1812; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1814 = 10'hf2 == _T_4[9:0] ? 8'h0 : _GEN_1813; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1815 = 10'hf3 == _T_4[9:0] ? 8'h0 : _GEN_1814; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1816 = 10'hf4 == _T_4[9:0] ? 8'hef : _GEN_1815; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1817 = 10'hf5 == _T_4[9:0] ? 8'hf0 : _GEN_1816; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1818 = 10'hf6 == _T_4[9:0] ? 8'h5f : _GEN_1817; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1819 = 10'hf7 == _T_4[9:0] ? 8'hf8 : _GEN_1818; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1820 = 10'hf8 == _T_4[9:0] ? 8'hef : _GEN_1819; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1821 = 10'hf9 == _T_4[9:0] ? 8'hf0 : _GEN_1820; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1822 = 10'hfa == _T_4[9:0] ? 8'h1f : _GEN_1821; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1823 = 10'hfb == _T_4[9:0] ? 8'hf5 : _GEN_1822; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1824 = 10'hfc == _T_4[9:0] ? 8'h93 : _GEN_1823; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1825 = 10'hfd == _T_4[9:0] ? 8'h7 : _GEN_1824; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1826 = 10'hfe == _T_4[9:0] ? 8'h5 : _GEN_1825; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1827 = 10'hff == _T_4[9:0] ? 8'h0 : _GEN_1826; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1828 = 10'h100 == _T_4[9:0] ? 8'he3 : _GEN_1827; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1829 = 10'h101 == _T_4[9:0] ? 8'h8c : _GEN_1828; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1830 = 10'h102 == _T_4[9:0] ? 8'h7 : _GEN_1829; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1831 = 10'h103 == _T_4[9:0] ? 8'hfe : _GEN_1830; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1832 = 10'h104 == _T_4[9:0] ? 8'hef : _GEN_1831; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1833 = 10'h105 == _T_4[9:0] ? 8'hf0 : _GEN_1832; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1834 = 10'h106 == _T_4[9:0] ? 8'h5f : _GEN_1833; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1835 = 10'h107 == _T_4[9:0] ? 8'hf1 : _GEN_1834; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1836 = 10'h108 == _T_4[9:0] ? 8'h93 : _GEN_1835; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1837 = 10'h109 == _T_4[9:0] ? 8'h7 : _GEN_1836; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1838 = 10'h10a == _T_4[9:0] ? 8'h5 : _GEN_1837; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1839 = 10'h10b == _T_4[9:0] ? 8'h0 : _GEN_1838; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1840 = 10'h10c == _T_4[9:0] ? 8'h13 : _GEN_1839; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1841 = 10'h10d == _T_4[9:0] ? 8'h85 : _GEN_1840; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1842 = 10'h10e == _T_4[9:0] ? 8'h7 : _GEN_1841; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1843 = 10'h10f == _T_4[9:0] ? 8'h0 : _GEN_1842; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1844 = 10'h110 == _T_4[9:0] ? 8'hef : _GEN_1843; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1845 = 10'h111 == _T_4[9:0] ? 8'hf0 : _GEN_1844; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1846 = 10'h112 == _T_4[9:0] ? 8'h9f : _GEN_1845; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1847 = 10'h113 == _T_4[9:0] ? 8'hf6 : _GEN_1846; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1848 = 10'h114 == _T_4[9:0] ? 8'h23 : _GEN_1847; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1849 = 10'h115 == _T_4[9:0] ? 8'h26 : _GEN_1848; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1850 = 10'h116 == _T_4[9:0] ? 8'h4 : _GEN_1849; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1851 = 10'h117 == _T_4[9:0] ? 8'hfe : _GEN_1850; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1852 = 10'h118 == _T_4[9:0] ? 8'h6f : _GEN_1851; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1853 = 10'h119 == _T_4[9:0] ? 8'h0 : _GEN_1852; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1854 = 10'h11a == _T_4[9:0] ? 8'h0 : _GEN_1853; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1855 = 10'h11b == _T_4[9:0] ? 8'h1 : _GEN_1854; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1856 = 10'h11c == _T_4[9:0] ? 8'h83 : _GEN_1855; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1857 = 10'h11d == _T_4[9:0] ? 8'h27 : _GEN_1856; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1858 = 10'h11e == _T_4[9:0] ? 8'hc4 : _GEN_1857; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1859 = 10'h11f == _T_4[9:0] ? 8'hfe : _GEN_1858; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1860 = 10'h120 == _T_4[9:0] ? 8'h93 : _GEN_1859; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1861 = 10'h121 == _T_4[9:0] ? 8'h87 : _GEN_1860; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1862 = 10'h122 == _T_4[9:0] ? 8'h17 : _GEN_1861; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1863 = 10'h123 == _T_4[9:0] ? 8'h0 : _GEN_1862; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1864 = 10'h124 == _T_4[9:0] ? 8'h23 : _GEN_1863; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1865 = 10'h125 == _T_4[9:0] ? 8'h26 : _GEN_1864; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1866 = 10'h126 == _T_4[9:0] ? 8'hf4 : _GEN_1865; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1867 = 10'h127 == _T_4[9:0] ? 8'hfe : _GEN_1866; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1868 = 10'h128 == _T_4[9:0] ? 8'h3 : _GEN_1867; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1869 = 10'h129 == _T_4[9:0] ? 8'h27 : _GEN_1868; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1870 = 10'h12a == _T_4[9:0] ? 8'hc4 : _GEN_1869; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1871 = 10'h12b == _T_4[9:0] ? 8'hfe : _GEN_1870; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1872 = 10'h12c == _T_4[9:0] ? 8'hb7 : _GEN_1871; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1873 = 10'h12d == _T_4[9:0] ? 8'h57 : _GEN_1872; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1874 = 10'h12e == _T_4[9:0] ? 8'h89 : _GEN_1873; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1875 = 10'h12f == _T_4[9:0] ? 8'h0 : _GEN_1874; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1876 = 10'h130 == _T_4[9:0] ? 8'h93 : _GEN_1875; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1877 = 10'h131 == _T_4[9:0] ? 8'h87 : _GEN_1876; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1878 = 10'h132 == _T_4[9:0] ? 8'hf7 : _GEN_1877; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1879 = 10'h133 == _T_4[9:0] ? 8'h43 : _GEN_1878; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1880 = 10'h134 == _T_4[9:0] ? 8'he3 : _GEN_1879; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1881 = 10'h135 == _T_4[9:0] ? 8'hd4 : _GEN_1880; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1882 = 10'h136 == _T_4[9:0] ? 8'he7 : _GEN_1881; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1883 = 10'h137 == _T_4[9:0] ? 8'hfe : _GEN_1882; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1884 = 10'h138 == _T_4[9:0] ? 8'h13 : _GEN_1883; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1885 = 10'h139 == _T_4[9:0] ? 8'h5 : _GEN_1884; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1886 = 10'h13a == _T_4[9:0] ? 8'h0 : _GEN_1885; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1887 = 10'h13b == _T_4[9:0] ? 8'h0 : _GEN_1886; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1888 = 10'h13c == _T_4[9:0] ? 8'hef : _GEN_1887; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1889 = 10'h13d == _T_4[9:0] ? 8'hf0 : _GEN_1888; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1890 = 10'h13e == _T_4[9:0] ? 8'hdf : _GEN_1889; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1891 = 10'h13f == _T_4[9:0] ? 8'hf3 : _GEN_1890; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1892 = 10'h140 == _T_4[9:0] ? 8'h6f : _GEN_1891; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1893 = 10'h141 == _T_4[9:0] ? 8'hf0 : _GEN_1892; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1894 = 10'h142 == _T_4[9:0] ? 8'h9f : _GEN_1893; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1895 = 10'h143 == _T_4[9:0] ? 8'hfb : _GEN_1894; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1896 = 10'h144 == _T_4[9:0] ? 8'h0 : _GEN_1895; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1897 = 10'h145 == _T_4[9:0] ? 8'h0 : _GEN_1896; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1898 = 10'h146 == _T_4[9:0] ? 8'h0 : _GEN_1897; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1899 = 10'h147 == _T_4[9:0] ? 8'h0 : _GEN_1898; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1900 = 10'h148 == _T_4[9:0] ? 8'h0 : _GEN_1899; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1901 = 10'h149 == _T_4[9:0] ? 8'h0 : _GEN_1900; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1902 = 10'h14a == _T_4[9:0] ? 8'h0 : _GEN_1901; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1903 = 10'h14b == _T_4[9:0] ? 8'h0 : _GEN_1902; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1904 = 10'h14c == _T_4[9:0] ? 8'h0 : _GEN_1903; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1905 = 10'h14d == _T_4[9:0] ? 8'h0 : _GEN_1904; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1906 = 10'h14e == _T_4[9:0] ? 8'h0 : _GEN_1905; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1907 = 10'h14f == _T_4[9:0] ? 8'h0 : _GEN_1906; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1908 = 10'h150 == _T_4[9:0] ? 8'h0 : _GEN_1907; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1909 = 10'h151 == _T_4[9:0] ? 8'h0 : _GEN_1908; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1910 = 10'h152 == _T_4[9:0] ? 8'h0 : _GEN_1909; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1911 = 10'h153 == _T_4[9:0] ? 8'h0 : _GEN_1910; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1912 = 10'h154 == _T_4[9:0] ? 8'h0 : _GEN_1911; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1913 = 10'h155 == _T_4[9:0] ? 8'h0 : _GEN_1912; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1914 = 10'h156 == _T_4[9:0] ? 8'h0 : _GEN_1913; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1915 = 10'h157 == _T_4[9:0] ? 8'h0 : _GEN_1914; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1916 = 10'h158 == _T_4[9:0] ? 8'h0 : _GEN_1915; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1917 = 10'h159 == _T_4[9:0] ? 8'h0 : _GEN_1916; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1918 = 10'h15a == _T_4[9:0] ? 8'h0 : _GEN_1917; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1919 = 10'h15b == _T_4[9:0] ? 8'h0 : _GEN_1918; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1920 = 10'h15c == _T_4[9:0] ? 8'h0 : _GEN_1919; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1921 = 10'h15d == _T_4[9:0] ? 8'h0 : _GEN_1920; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1922 = 10'h15e == _T_4[9:0] ? 8'h0 : _GEN_1921; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1923 = 10'h15f == _T_4[9:0] ? 8'h0 : _GEN_1922; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1924 = 10'h160 == _T_4[9:0] ? 8'h0 : _GEN_1923; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1925 = 10'h161 == _T_4[9:0] ? 8'h0 : _GEN_1924; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1926 = 10'h162 == _T_4[9:0] ? 8'h0 : _GEN_1925; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1927 = 10'h163 == _T_4[9:0] ? 8'h0 : _GEN_1926; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1928 = 10'h164 == _T_4[9:0] ? 8'h0 : _GEN_1927; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1929 = 10'h165 == _T_4[9:0] ? 8'h0 : _GEN_1928; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1930 = 10'h166 == _T_4[9:0] ? 8'h0 : _GEN_1929; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1931 = 10'h167 == _T_4[9:0] ? 8'h0 : _GEN_1930; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1932 = 10'h168 == _T_4[9:0] ? 8'h0 : _GEN_1931; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1933 = 10'h169 == _T_4[9:0] ? 8'h0 : _GEN_1932; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1934 = 10'h16a == _T_4[9:0] ? 8'h0 : _GEN_1933; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1935 = 10'h16b == _T_4[9:0] ? 8'h0 : _GEN_1934; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1936 = 10'h16c == _T_4[9:0] ? 8'h0 : _GEN_1935; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1937 = 10'h16d == _T_4[9:0] ? 8'h0 : _GEN_1936; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1938 = 10'h16e == _T_4[9:0] ? 8'h0 : _GEN_1937; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1939 = 10'h16f == _T_4[9:0] ? 8'h0 : _GEN_1938; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1940 = 10'h170 == _T_4[9:0] ? 8'h0 : _GEN_1939; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1941 = 10'h171 == _T_4[9:0] ? 8'h0 : _GEN_1940; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1942 = 10'h172 == _T_4[9:0] ? 8'h0 : _GEN_1941; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1943 = 10'h173 == _T_4[9:0] ? 8'h0 : _GEN_1942; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1944 = 10'h174 == _T_4[9:0] ? 8'h0 : _GEN_1943; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1945 = 10'h175 == _T_4[9:0] ? 8'h0 : _GEN_1944; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1946 = 10'h176 == _T_4[9:0] ? 8'h0 : _GEN_1945; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1947 = 10'h177 == _T_4[9:0] ? 8'h0 : _GEN_1946; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1948 = 10'h178 == _T_4[9:0] ? 8'h0 : _GEN_1947; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1949 = 10'h179 == _T_4[9:0] ? 8'h0 : _GEN_1948; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1950 = 10'h17a == _T_4[9:0] ? 8'h0 : _GEN_1949; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1951 = 10'h17b == _T_4[9:0] ? 8'h0 : _GEN_1950; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1952 = 10'h17c == _T_4[9:0] ? 8'h0 : _GEN_1951; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1953 = 10'h17d == _T_4[9:0] ? 8'h0 : _GEN_1952; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1954 = 10'h17e == _T_4[9:0] ? 8'h0 : _GEN_1953; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1955 = 10'h17f == _T_4[9:0] ? 8'h0 : _GEN_1954; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1956 = 10'h180 == _T_4[9:0] ? 8'h0 : _GEN_1955; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1957 = 10'h181 == _T_4[9:0] ? 8'h0 : _GEN_1956; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1958 = 10'h182 == _T_4[9:0] ? 8'h0 : _GEN_1957; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1959 = 10'h183 == _T_4[9:0] ? 8'h0 : _GEN_1958; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1960 = 10'h184 == _T_4[9:0] ? 8'h0 : _GEN_1959; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1961 = 10'h185 == _T_4[9:0] ? 8'h0 : _GEN_1960; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1962 = 10'h186 == _T_4[9:0] ? 8'h0 : _GEN_1961; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1963 = 10'h187 == _T_4[9:0] ? 8'h0 : _GEN_1962; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1964 = 10'h188 == _T_4[9:0] ? 8'h0 : _GEN_1963; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1965 = 10'h189 == _T_4[9:0] ? 8'h0 : _GEN_1964; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1966 = 10'h18a == _T_4[9:0] ? 8'h0 : _GEN_1965; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1967 = 10'h18b == _T_4[9:0] ? 8'h0 : _GEN_1966; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1968 = 10'h18c == _T_4[9:0] ? 8'h0 : _GEN_1967; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1969 = 10'h18d == _T_4[9:0] ? 8'h0 : _GEN_1968; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1970 = 10'h18e == _T_4[9:0] ? 8'h0 : _GEN_1969; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1971 = 10'h18f == _T_4[9:0] ? 8'h0 : _GEN_1970; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1972 = 10'h190 == _T_4[9:0] ? 8'h0 : _GEN_1971; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1973 = 10'h191 == _T_4[9:0] ? 8'h0 : _GEN_1972; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1974 = 10'h192 == _T_4[9:0] ? 8'h0 : _GEN_1973; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1975 = 10'h193 == _T_4[9:0] ? 8'h0 : _GEN_1974; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1976 = 10'h194 == _T_4[9:0] ? 8'h0 : _GEN_1975; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1977 = 10'h195 == _T_4[9:0] ? 8'h0 : _GEN_1976; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1978 = 10'h196 == _T_4[9:0] ? 8'h0 : _GEN_1977; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1979 = 10'h197 == _T_4[9:0] ? 8'h0 : _GEN_1978; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1980 = 10'h198 == _T_4[9:0] ? 8'h0 : _GEN_1979; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1981 = 10'h199 == _T_4[9:0] ? 8'h0 : _GEN_1980; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1982 = 10'h19a == _T_4[9:0] ? 8'h0 : _GEN_1981; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1983 = 10'h19b == _T_4[9:0] ? 8'h0 : _GEN_1982; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1984 = 10'h19c == _T_4[9:0] ? 8'h0 : _GEN_1983; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1985 = 10'h19d == _T_4[9:0] ? 8'h0 : _GEN_1984; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1986 = 10'h19e == _T_4[9:0] ? 8'h0 : _GEN_1985; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1987 = 10'h19f == _T_4[9:0] ? 8'h0 : _GEN_1986; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1988 = 10'h1a0 == _T_4[9:0] ? 8'h0 : _GEN_1987; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1989 = 10'h1a1 == _T_4[9:0] ? 8'h0 : _GEN_1988; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1990 = 10'h1a2 == _T_4[9:0] ? 8'h0 : _GEN_1989; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1991 = 10'h1a3 == _T_4[9:0] ? 8'h0 : _GEN_1990; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1992 = 10'h1a4 == _T_4[9:0] ? 8'h0 : _GEN_1991; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1993 = 10'h1a5 == _T_4[9:0] ? 8'h0 : _GEN_1992; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1994 = 10'h1a6 == _T_4[9:0] ? 8'h0 : _GEN_1993; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1995 = 10'h1a7 == _T_4[9:0] ? 8'h0 : _GEN_1994; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1996 = 10'h1a8 == _T_4[9:0] ? 8'h0 : _GEN_1995; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1997 = 10'h1a9 == _T_4[9:0] ? 8'h0 : _GEN_1996; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1998 = 10'h1aa == _T_4[9:0] ? 8'h0 : _GEN_1997; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1999 = 10'h1ab == _T_4[9:0] ? 8'h0 : _GEN_1998; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2000 = 10'h1ac == _T_4[9:0] ? 8'h0 : _GEN_1999; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2001 = 10'h1ad == _T_4[9:0] ? 8'h0 : _GEN_2000; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2002 = 10'h1ae == _T_4[9:0] ? 8'h0 : _GEN_2001; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2003 = 10'h1af == _T_4[9:0] ? 8'h0 : _GEN_2002; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2004 = 10'h1b0 == _T_4[9:0] ? 8'h0 : _GEN_2003; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2005 = 10'h1b1 == _T_4[9:0] ? 8'h0 : _GEN_2004; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2006 = 10'h1b2 == _T_4[9:0] ? 8'h0 : _GEN_2005; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2007 = 10'h1b3 == _T_4[9:0] ? 8'h0 : _GEN_2006; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2008 = 10'h1b4 == _T_4[9:0] ? 8'h0 : _GEN_2007; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2009 = 10'h1b5 == _T_4[9:0] ? 8'h0 : _GEN_2008; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2010 = 10'h1b6 == _T_4[9:0] ? 8'h0 : _GEN_2009; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2011 = 10'h1b7 == _T_4[9:0] ? 8'h0 : _GEN_2010; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2012 = 10'h1b8 == _T_4[9:0] ? 8'h0 : _GEN_2011; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2013 = 10'h1b9 == _T_4[9:0] ? 8'h0 : _GEN_2012; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2014 = 10'h1ba == _T_4[9:0] ? 8'h0 : _GEN_2013; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2015 = 10'h1bb == _T_4[9:0] ? 8'h0 : _GEN_2014; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2016 = 10'h1bc == _T_4[9:0] ? 8'h0 : _GEN_2015; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2017 = 10'h1bd == _T_4[9:0] ? 8'h0 : _GEN_2016; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2018 = 10'h1be == _T_4[9:0] ? 8'h0 : _GEN_2017; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2019 = 10'h1bf == _T_4[9:0] ? 8'h0 : _GEN_2018; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2020 = 10'h1c0 == _T_4[9:0] ? 8'h0 : _GEN_2019; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2021 = 10'h1c1 == _T_4[9:0] ? 8'h0 : _GEN_2020; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2022 = 10'h1c2 == _T_4[9:0] ? 8'h0 : _GEN_2021; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2023 = 10'h1c3 == _T_4[9:0] ? 8'h0 : _GEN_2022; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2024 = 10'h1c4 == _T_4[9:0] ? 8'h0 : _GEN_2023; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2025 = 10'h1c5 == _T_4[9:0] ? 8'h0 : _GEN_2024; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2026 = 10'h1c6 == _T_4[9:0] ? 8'h0 : _GEN_2025; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2027 = 10'h1c7 == _T_4[9:0] ? 8'h0 : _GEN_2026; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2028 = 10'h1c8 == _T_4[9:0] ? 8'h0 : _GEN_2027; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2029 = 10'h1c9 == _T_4[9:0] ? 8'h0 : _GEN_2028; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2030 = 10'h1ca == _T_4[9:0] ? 8'h0 : _GEN_2029; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2031 = 10'h1cb == _T_4[9:0] ? 8'h0 : _GEN_2030; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2032 = 10'h1cc == _T_4[9:0] ? 8'h0 : _GEN_2031; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2033 = 10'h1cd == _T_4[9:0] ? 8'h0 : _GEN_2032; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2034 = 10'h1ce == _T_4[9:0] ? 8'h0 : _GEN_2033; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2035 = 10'h1cf == _T_4[9:0] ? 8'h0 : _GEN_2034; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2036 = 10'h1d0 == _T_4[9:0] ? 8'h0 : _GEN_2035; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2037 = 10'h1d1 == _T_4[9:0] ? 8'h0 : _GEN_2036; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2038 = 10'h1d2 == _T_4[9:0] ? 8'h0 : _GEN_2037; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2039 = 10'h1d3 == _T_4[9:0] ? 8'h0 : _GEN_2038; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2040 = 10'h1d4 == _T_4[9:0] ? 8'h0 : _GEN_2039; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2041 = 10'h1d5 == _T_4[9:0] ? 8'h0 : _GEN_2040; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2042 = 10'h1d6 == _T_4[9:0] ? 8'h0 : _GEN_2041; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2043 = 10'h1d7 == _T_4[9:0] ? 8'h0 : _GEN_2042; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2044 = 10'h1d8 == _T_4[9:0] ? 8'h0 : _GEN_2043; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2045 = 10'h1d9 == _T_4[9:0] ? 8'h0 : _GEN_2044; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2046 = 10'h1da == _T_4[9:0] ? 8'h0 : _GEN_2045; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2047 = 10'h1db == _T_4[9:0] ? 8'h0 : _GEN_2046; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2048 = 10'h1dc == _T_4[9:0] ? 8'h0 : _GEN_2047; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2049 = 10'h1dd == _T_4[9:0] ? 8'h0 : _GEN_2048; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2050 = 10'h1de == _T_4[9:0] ? 8'h0 : _GEN_2049; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2051 = 10'h1df == _T_4[9:0] ? 8'h0 : _GEN_2050; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2052 = 10'h1e0 == _T_4[9:0] ? 8'h0 : _GEN_2051; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2053 = 10'h1e1 == _T_4[9:0] ? 8'h0 : _GEN_2052; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2054 = 10'h1e2 == _T_4[9:0] ? 8'h0 : _GEN_2053; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2055 = 10'h1e3 == _T_4[9:0] ? 8'h0 : _GEN_2054; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2056 = 10'h1e4 == _T_4[9:0] ? 8'h0 : _GEN_2055; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2057 = 10'h1e5 == _T_4[9:0] ? 8'h0 : _GEN_2056; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2058 = 10'h1e6 == _T_4[9:0] ? 8'h0 : _GEN_2057; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2059 = 10'h1e7 == _T_4[9:0] ? 8'h0 : _GEN_2058; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2060 = 10'h1e8 == _T_4[9:0] ? 8'h0 : _GEN_2059; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2061 = 10'h1e9 == _T_4[9:0] ? 8'h0 : _GEN_2060; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2062 = 10'h1ea == _T_4[9:0] ? 8'h0 : _GEN_2061; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2063 = 10'h1eb == _T_4[9:0] ? 8'h0 : _GEN_2062; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2064 = 10'h1ec == _T_4[9:0] ? 8'h0 : _GEN_2063; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2065 = 10'h1ed == _T_4[9:0] ? 8'h0 : _GEN_2064; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2066 = 10'h1ee == _T_4[9:0] ? 8'h0 : _GEN_2065; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2067 = 10'h1ef == _T_4[9:0] ? 8'h0 : _GEN_2066; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2068 = 10'h1f0 == _T_4[9:0] ? 8'h0 : _GEN_2067; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2069 = 10'h1f1 == _T_4[9:0] ? 8'h0 : _GEN_2068; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2070 = 10'h1f2 == _T_4[9:0] ? 8'h0 : _GEN_2069; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2071 = 10'h1f3 == _T_4[9:0] ? 8'h0 : _GEN_2070; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2072 = 10'h1f4 == _T_4[9:0] ? 8'h0 : _GEN_2071; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2073 = 10'h1f5 == _T_4[9:0] ? 8'h0 : _GEN_2072; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2074 = 10'h1f6 == _T_4[9:0] ? 8'h0 : _GEN_2073; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2075 = 10'h1f7 == _T_4[9:0] ? 8'h0 : _GEN_2074; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2076 = 10'h1f8 == _T_4[9:0] ? 8'h0 : _GEN_2075; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2077 = 10'h1f9 == _T_4[9:0] ? 8'h0 : _GEN_2076; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2078 = 10'h1fa == _T_4[9:0] ? 8'h0 : _GEN_2077; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2079 = 10'h1fb == _T_4[9:0] ? 8'h0 : _GEN_2078; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2080 = 10'h1fc == _T_4[9:0] ? 8'h0 : _GEN_2079; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2081 = 10'h1fd == _T_4[9:0] ? 8'h0 : _GEN_2080; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2082 = 10'h1fe == _T_4[9:0] ? 8'h0 : _GEN_2081; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2083 = 10'h1ff == _T_4[9:0] ? 8'h0 : _GEN_2082; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2084 = 10'h200 == _T_4[9:0] ? 8'h0 : _GEN_2083; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2085 = 10'h201 == _T_4[9:0] ? 8'h0 : _GEN_2084; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2086 = 10'h202 == _T_4[9:0] ? 8'h0 : _GEN_2085; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2087 = 10'h203 == _T_4[9:0] ? 8'h0 : _GEN_2086; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2088 = 10'h204 == _T_4[9:0] ? 8'h0 : _GEN_2087; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2089 = 10'h205 == _T_4[9:0] ? 8'h0 : _GEN_2088; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2090 = 10'h206 == _T_4[9:0] ? 8'h0 : _GEN_2089; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2091 = 10'h207 == _T_4[9:0] ? 8'h0 : _GEN_2090; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2092 = 10'h208 == _T_4[9:0] ? 8'h0 : _GEN_2091; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2093 = 10'h209 == _T_4[9:0] ? 8'h0 : _GEN_2092; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2094 = 10'h20a == _T_4[9:0] ? 8'h0 : _GEN_2093; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2095 = 10'h20b == _T_4[9:0] ? 8'h0 : _GEN_2094; // @[Cat.scala 29:58]
  wire [31:0] _T_16 = pc + 32'h4; // @[IF.scala 47:14]
  assign out_pc = pc; // @[IF.scala 42:10]
  assign out_instr = {_GEN_1571,_GEN_2095,_GEN_523,_GEN_1047}; // @[IF.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h0;
    end else if (ctrl_pcEn) begin
      if (in_branch) begin
        pc <= in_pcNext;
      end else begin
        pc <= _T_16;
      end
    end
  end
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_registerS1Index,
  input  [4:0]  io_registerS2Index,
  input  [4:0]  io_registerWIndex,
  input  [31:0] io_registerWData,
  input         io_writeEn,
  output [31:0] io_registerS1Data,
  output [31:0] io_registerS2Data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regFile_1; // @[RegFile.scala 20:24]
  reg [31:0] regFile_2; // @[RegFile.scala 20:24]
  reg [31:0] regFile_3; // @[RegFile.scala 20:24]
  reg [31:0] regFile_4; // @[RegFile.scala 20:24]
  reg [31:0] regFile_5; // @[RegFile.scala 20:24]
  reg [31:0] regFile_6; // @[RegFile.scala 20:24]
  reg [31:0] regFile_7; // @[RegFile.scala 20:24]
  reg [31:0] regFile_8; // @[RegFile.scala 20:24]
  reg [31:0] regFile_9; // @[RegFile.scala 20:24]
  reg [31:0] regFile_10; // @[RegFile.scala 20:24]
  reg [31:0] regFile_11; // @[RegFile.scala 20:24]
  reg [31:0] regFile_12; // @[RegFile.scala 20:24]
  reg [31:0] regFile_13; // @[RegFile.scala 20:24]
  reg [31:0] regFile_14; // @[RegFile.scala 20:24]
  reg [31:0] regFile_15; // @[RegFile.scala 20:24]
  reg [31:0] regFile_16; // @[RegFile.scala 20:24]
  reg [31:0] regFile_17; // @[RegFile.scala 20:24]
  reg [31:0] regFile_18; // @[RegFile.scala 20:24]
  reg [31:0] regFile_19; // @[RegFile.scala 20:24]
  reg [31:0] regFile_20; // @[RegFile.scala 20:24]
  reg [31:0] regFile_21; // @[RegFile.scala 20:24]
  reg [31:0] regFile_22; // @[RegFile.scala 20:24]
  reg [31:0] regFile_23; // @[RegFile.scala 20:24]
  reg [31:0] regFile_24; // @[RegFile.scala 20:24]
  reg [31:0] regFile_25; // @[RegFile.scala 20:24]
  reg [31:0] regFile_26; // @[RegFile.scala 20:24]
  reg [31:0] regFile_27; // @[RegFile.scala 20:24]
  reg [31:0] regFile_28; // @[RegFile.scala 20:24]
  reg [31:0] regFile_29; // @[RegFile.scala 20:24]
  reg [31:0] regFile_30; // @[RegFile.scala 20:24]
  reg [31:0] regFile_31; // @[RegFile.scala 20:24]
  wire [31:0] _GEN_65 = 5'h1 == io_registerS1Index ? $signed(regFile_1) : $signed(32'sh0); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_66 = 5'h2 == io_registerS1Index ? $signed(regFile_2) : $signed(_GEN_65); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_67 = 5'h3 == io_registerS1Index ? $signed(regFile_3) : $signed(_GEN_66); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_68 = 5'h4 == io_registerS1Index ? $signed(regFile_4) : $signed(_GEN_67); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_69 = 5'h5 == io_registerS1Index ? $signed(regFile_5) : $signed(_GEN_68); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_70 = 5'h6 == io_registerS1Index ? $signed(regFile_6) : $signed(_GEN_69); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_71 = 5'h7 == io_registerS1Index ? $signed(regFile_7) : $signed(_GEN_70); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_72 = 5'h8 == io_registerS1Index ? $signed(regFile_8) : $signed(_GEN_71); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_73 = 5'h9 == io_registerS1Index ? $signed(regFile_9) : $signed(_GEN_72); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_74 = 5'ha == io_registerS1Index ? $signed(regFile_10) : $signed(_GEN_73); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_75 = 5'hb == io_registerS1Index ? $signed(regFile_11) : $signed(_GEN_74); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_76 = 5'hc == io_registerS1Index ? $signed(regFile_12) : $signed(_GEN_75); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_77 = 5'hd == io_registerS1Index ? $signed(regFile_13) : $signed(_GEN_76); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_78 = 5'he == io_registerS1Index ? $signed(regFile_14) : $signed(_GEN_77); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_79 = 5'hf == io_registerS1Index ? $signed(regFile_15) : $signed(_GEN_78); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_80 = 5'h10 == io_registerS1Index ? $signed(regFile_16) : $signed(_GEN_79); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_81 = 5'h11 == io_registerS1Index ? $signed(regFile_17) : $signed(_GEN_80); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_82 = 5'h12 == io_registerS1Index ? $signed(regFile_18) : $signed(_GEN_81); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_83 = 5'h13 == io_registerS1Index ? $signed(regFile_19) : $signed(_GEN_82); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_84 = 5'h14 == io_registerS1Index ? $signed(regFile_20) : $signed(_GEN_83); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_85 = 5'h15 == io_registerS1Index ? $signed(regFile_21) : $signed(_GEN_84); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_86 = 5'h16 == io_registerS1Index ? $signed(regFile_22) : $signed(_GEN_85); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_87 = 5'h17 == io_registerS1Index ? $signed(regFile_23) : $signed(_GEN_86); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_88 = 5'h18 == io_registerS1Index ? $signed(regFile_24) : $signed(_GEN_87); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_89 = 5'h19 == io_registerS1Index ? $signed(regFile_25) : $signed(_GEN_88); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_90 = 5'h1a == io_registerS1Index ? $signed(regFile_26) : $signed(_GEN_89); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_91 = 5'h1b == io_registerS1Index ? $signed(regFile_27) : $signed(_GEN_90); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_92 = 5'h1c == io_registerS1Index ? $signed(regFile_28) : $signed(_GEN_91); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_93 = 5'h1d == io_registerS1Index ? $signed(regFile_29) : $signed(_GEN_92); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_94 = 5'h1e == io_registerS1Index ? $signed(regFile_30) : $signed(_GEN_93); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_95 = 5'h1f == io_registerS1Index ? $signed(regFile_31) : $signed(_GEN_94); // @[RegFile.scala 27:21]
  wire [31:0] _GEN_97 = 5'h1 == io_registerS2Index ? $signed(regFile_1) : $signed(32'sh0); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_98 = 5'h2 == io_registerS2Index ? $signed(regFile_2) : $signed(_GEN_97); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_99 = 5'h3 == io_registerS2Index ? $signed(regFile_3) : $signed(_GEN_98); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_100 = 5'h4 == io_registerS2Index ? $signed(regFile_4) : $signed(_GEN_99); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_101 = 5'h5 == io_registerS2Index ? $signed(regFile_5) : $signed(_GEN_100); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_102 = 5'h6 == io_registerS2Index ? $signed(regFile_6) : $signed(_GEN_101); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_103 = 5'h7 == io_registerS2Index ? $signed(regFile_7) : $signed(_GEN_102); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_104 = 5'h8 == io_registerS2Index ? $signed(regFile_8) : $signed(_GEN_103); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_105 = 5'h9 == io_registerS2Index ? $signed(regFile_9) : $signed(_GEN_104); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_106 = 5'ha == io_registerS2Index ? $signed(regFile_10) : $signed(_GEN_105); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_107 = 5'hb == io_registerS2Index ? $signed(regFile_11) : $signed(_GEN_106); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_108 = 5'hc == io_registerS2Index ? $signed(regFile_12) : $signed(_GEN_107); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_109 = 5'hd == io_registerS2Index ? $signed(regFile_13) : $signed(_GEN_108); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_110 = 5'he == io_registerS2Index ? $signed(regFile_14) : $signed(_GEN_109); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_111 = 5'hf == io_registerS2Index ? $signed(regFile_15) : $signed(_GEN_110); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_112 = 5'h10 == io_registerS2Index ? $signed(regFile_16) : $signed(_GEN_111); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_113 = 5'h11 == io_registerS2Index ? $signed(regFile_17) : $signed(_GEN_112); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_114 = 5'h12 == io_registerS2Index ? $signed(regFile_18) : $signed(_GEN_113); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_115 = 5'h13 == io_registerS2Index ? $signed(regFile_19) : $signed(_GEN_114); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_116 = 5'h14 == io_registerS2Index ? $signed(regFile_20) : $signed(_GEN_115); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_117 = 5'h15 == io_registerS2Index ? $signed(regFile_21) : $signed(_GEN_116); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_118 = 5'h16 == io_registerS2Index ? $signed(regFile_22) : $signed(_GEN_117); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_119 = 5'h17 == io_registerS2Index ? $signed(regFile_23) : $signed(_GEN_118); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_120 = 5'h18 == io_registerS2Index ? $signed(regFile_24) : $signed(_GEN_119); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_121 = 5'h19 == io_registerS2Index ? $signed(regFile_25) : $signed(_GEN_120); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_122 = 5'h1a == io_registerS2Index ? $signed(regFile_26) : $signed(_GEN_121); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_123 = 5'h1b == io_registerS2Index ? $signed(regFile_27) : $signed(_GEN_122); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_124 = 5'h1c == io_registerS2Index ? $signed(regFile_28) : $signed(_GEN_123); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_125 = 5'h1d == io_registerS2Index ? $signed(regFile_29) : $signed(_GEN_124); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_126 = 5'h1e == io_registerS2Index ? $signed(regFile_30) : $signed(_GEN_125); // @[RegFile.scala 28:21]
  wire [31:0] _GEN_127 = 5'h1f == io_registerS2Index ? $signed(regFile_31) : $signed(_GEN_126); // @[RegFile.scala 28:21]
  wire  _T_1 = io_registerS1Index == io_registerWIndex; // @[RegFile.scala 30:27]
  wire  _T_2 = io_registerS1Index != 5'h0; // @[RegFile.scala 30:71]
  wire  _T_3 = _T_1 & _T_2; // @[RegFile.scala 30:49]
  wire  _T_4 = _T_3 & io_writeEn; // @[RegFile.scala 30:79]
  wire  _T_5 = io_registerS2Index == io_registerWIndex; // @[RegFile.scala 33:27]
  wire  _T_6 = io_registerS2Index != 5'h0; // @[RegFile.scala 33:71]
  wire  _T_7 = _T_5 & _T_6; // @[RegFile.scala 33:49]
  wire  _T_8 = _T_7 & io_writeEn; // @[RegFile.scala 33:79]
  assign io_registerS1Data = _T_4 ? $signed(io_registerWData) : $signed(_GEN_95); // @[RegFile.scala 27:21 RegFile.scala 31:23]
  assign io_registerS2Data = _T_8 ? $signed(io_registerWData) : $signed(_GEN_127); // @[RegFile.scala 28:21 RegFile.scala 34:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regFile_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regFile_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regFile_3 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regFile_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regFile_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regFile_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regFile_7 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regFile_8 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regFile_9 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regFile_10 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regFile_11 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regFile_12 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regFile_13 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regFile_14 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regFile_15 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regFile_16 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regFile_17 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regFile_18 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regFile_19 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regFile_20 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regFile_21 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regFile_22 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regFile_23 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regFile_24 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regFile_25 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regFile_26 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regFile_27 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regFile_28 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regFile_29 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regFile_30 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regFile_31 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regFile_1 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1 == io_registerWIndex) begin
        regFile_1 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_2 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h2 == io_registerWIndex) begin
        regFile_2 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_3 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h3 == io_registerWIndex) begin
        regFile_3 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_4 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h4 == io_registerWIndex) begin
        regFile_4 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_5 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h5 == io_registerWIndex) begin
        regFile_5 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_6 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h6 == io_registerWIndex) begin
        regFile_6 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_7 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h7 == io_registerWIndex) begin
        regFile_7 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_8 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h8 == io_registerWIndex) begin
        regFile_8 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_9 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h9 == io_registerWIndex) begin
        regFile_9 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_10 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'ha == io_registerWIndex) begin
        regFile_10 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_11 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hb == io_registerWIndex) begin
        regFile_11 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_12 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hc == io_registerWIndex) begin
        regFile_12 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_13 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hd == io_registerWIndex) begin
        regFile_13 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_14 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'he == io_registerWIndex) begin
        regFile_14 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_15 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hf == io_registerWIndex) begin
        regFile_15 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_16 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h10 == io_registerWIndex) begin
        regFile_16 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_17 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h11 == io_registerWIndex) begin
        regFile_17 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_18 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h12 == io_registerWIndex) begin
        regFile_18 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_19 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h13 == io_registerWIndex) begin
        regFile_19 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_20 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h14 == io_registerWIndex) begin
        regFile_20 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_21 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h15 == io_registerWIndex) begin
        regFile_21 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_22 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h16 == io_registerWIndex) begin
        regFile_22 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_23 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h17 == io_registerWIndex) begin
        regFile_23 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_24 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h18 == io_registerWIndex) begin
        regFile_24 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_25 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h19 == io_registerWIndex) begin
        regFile_25 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_26 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1a == io_registerWIndex) begin
        regFile_26 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_27 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1b == io_registerWIndex) begin
        regFile_27 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_28 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1c == io_registerWIndex) begin
        regFile_28 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_29 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1d == io_registerWIndex) begin
        regFile_29 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_30 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1e == io_registerWIndex) begin
        regFile_30 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_31 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1f == io_registerWIndex) begin
        regFile_31 <= io_registerWData;
      end
    end
  end
endmodule
module ImmGen(
  input  [31:0] io_instruction,
  output [31:0] io_immediate
);
  wire [2:0] funct3 = io_instruction[14:12]; // @[ImmGen.scala 13:30]
  wire [11:0] Itype = io_instruction[31:20]; // @[ImmGen.scala 19:29]
  wire [9:0] _T_45 = {io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31]}; // @[ImmGen.scala 21:71]
  wire [31:0] _T_57 = {_T_45,_T_45,Itype}; // @[ImmGen.scala 21:88]
  wire  _T_58 = funct3 == 3'h2; // @[ImmGen.scala 22:15]
  wire  _T_59 = funct3 == 3'h3; // @[ImmGen.scala 22:33]
  wire  _T_60 = _T_58 | _T_59; // @[ImmGen.scala 22:23]
  wire [11:0] _T_61 = io_instruction[31:20]; // @[ImmGen.scala 23:33]
  wire [31:0] _GEN_0 = _T_60 ? $signed({{20{_T_61[11]}},_T_61}) : $signed(_T_57); // @[ImmGen.scala 22:42]
  wire  _T_63 = 7'h37 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [31:0] _T_64 = {io_instruction[31:12],12'h0}; // @[ImmGen.scala 29:35]
  wire  _T_65 = 7'h17 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_67 = 7'h6f == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [30:0] _T_90 = {_T_45,io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:22],2'h0}; // @[ImmGen.scala 35:103]
  wire  _T_91 = 7'h23 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [31:0] _T_133 = {_T_45,_T_45,io_instruction[31:25],io_instruction[11:7]}; // @[ImmGen.scala 38:92]
  wire  _T_134 = 7'h63 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [8:0] _T_161 = {io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31]}; // @[ImmGen.scala 41:75]
  wire [17:0] _T_170 = {io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],_T_161}; // @[ImmGen.scala 41:75]
  wire [30:0] _T_173 = {_T_170,io_instruction[31],io_instruction[7],io_instruction[30:25],io_instruction[11:8],1'h0}; // @[ImmGen.scala 41:103]
  wire [31:0] _GEN_1 = _T_134 ? $signed({{1{_T_173[30]}},_T_173}) : $signed(_GEN_0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_91 ? $signed(_T_133) : $signed(_GEN_1); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_3 = _T_67 ? $signed({{1{_T_90[30]}},_T_90}) : $signed(_GEN_2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_4 = _T_65 ? $signed(_T_64) : $signed(_GEN_3); // @[Conditional.scala 39:67]
  assign io_immediate = _T_63 ? $signed(_T_64) : $signed(_GEN_4); // @[ImmGen.scala 21:16 ImmGen.scala 23:18 ImmGen.scala 29:20 ImmGen.scala 32:20 ImmGen.scala 35:20 ImmGen.scala 38:20 ImmGen.scala 41:20]
endmodule
module ID(
  input         clock,
  input         reset,
  input  [31:0] in_pc,
  input  [31:0] in_instr,
  output [31:0] out_pc,
  output [31:0] out_imm,
  output [31:0] out_regOp1,
  output [31:0] out_regOp2,
  output [4:0]  out_rs1,
  output [4:0]  out_rs2,
  output [4:0]  out_rd,
  output [3:0]  out_aluOp,
  output [1:0]  out_aluSrc1,
  output [1:0]  out_aluSrc2,
  output        out_brSrc,
  output        out_pcSrc,
  output        out_wb,
  output        out_wbSrc,
  output [3:0]  out_mem,
  output        out_jump,
  output [2:0]  out_funct3,
  input  [4:0]  wb_rd,
  input  [31:0] wb_res,
  input         wb_wb,
  input         ctrl_flushID,
  output [31:0] ctrl_instr
);
  wire  regFile_clock; // @[ID.scala 21:23]
  wire  regFile_reset; // @[ID.scala 21:23]
  wire [4:0] regFile_io_registerS1Index; // @[ID.scala 21:23]
  wire [4:0] regFile_io_registerS2Index; // @[ID.scala 21:23]
  wire [4:0] regFile_io_registerWIndex; // @[ID.scala 21:23]
  wire [31:0] regFile_io_registerWData; // @[ID.scala 21:23]
  wire  regFile_io_writeEn; // @[ID.scala 21:23]
  wire [31:0] regFile_io_registerS1Data; // @[ID.scala 21:23]
  wire [31:0] regFile_io_registerS2Data; // @[ID.scala 21:23]
  wire [31:0] immGen_io_instruction; // @[ID.scala 23:22]
  wire [31:0] immGen_io_immediate; // @[ID.scala 23:22]
  wire [6:0] opcode = in_instr[6:0]; // @[ID.scala 25:24]
  wire [2:0] funct3 = in_instr[14:12]; // @[ID.scala 26:24]
  wire  _T_1 = 7'h3 == opcode; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h0 == funct3; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h4 == funct3; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h1 == funct3; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h5 == funct3; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h2 == funct3; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_0 = _T_6 ? 3'h7 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1 = _T_5 ? 3'h2 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_4 ? 3'h6 : _GEN_1; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_3 = _T_3 ? 3'h1 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_2 ? 3'h5 : _GEN_3; // @[Conditional.scala 40:58]
  wire  _T_7 = 7'h23 == opcode; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_5 = _T_6 ? 4'hb : 4'h0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_6 = _T_4 ? 4'ha : _GEN_5; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_7 = _T_2 ? 4'h9 : _GEN_6; // @[Conditional.scala 40:58]
  wire  _T_11 = 7'h13 == opcode; // @[Conditional.scala 37:30]
  wire  _T_15 = 3'h3 == funct3; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_8 = in_instr[30] ? 4'h4 : 4'h3; // @[ID.scala 118:30]
  wire  _T_19 = 3'h6 == funct3; // @[Conditional.scala 37:30]
  wire  _T_20 = 3'h7 == funct3; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_9 = _T_20 ? 4'h5 : 4'h0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_10 = _T_19 ? 4'h6 : _GEN_9; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_11 = _T_5 ? _GEN_8 : _GEN_10; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_12 = _T_3 ? 4'h7 : _GEN_11; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_13 = _T_15 ? 4'h8 : _GEN_12; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_14 = _T_6 ? 4'h8 : _GEN_13; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_15 = _T_4 ? 4'h2 : _GEN_14; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_16 = _T_2 ? 4'h0 : _GEN_15; // @[Conditional.scala 40:58]
  wire  _T_21 = 7'h33 == opcode; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_17 = in_instr[30] ? 4'h1 : 4'h0; // @[ID.scala 135:30]
  wire [3:0] _GEN_26 = _T_2 ? _GEN_17 : _GEN_15; // @[Conditional.scala 40:58]
  wire  _T_32 = 7'h17 == opcode; // @[Conditional.scala 37:30]
  wire  _T_33 = 7'h37 == opcode; // @[Conditional.scala 37:30]
  wire  _T_34 = 7'h63 == opcode; // @[Conditional.scala 37:30]
  wire  _T_35 = 7'h6f == opcode; // @[Conditional.scala 37:30]
  wire  _T_36 = 7'h67 == opcode; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_28 = _T_36 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_35 | _T_36; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_30 = _T_35 ? 2'h1 : _GEN_28; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_31 = _T_35 ? 2'h2 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_32 = _T_35 ? 1'h0 : _T_36; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_34 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_34 | _GEN_29; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_35 = _T_34 ? 2'h0 : _GEN_30; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_36 = _T_34 ? 2'h0 : _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_34 ? 1'h0 : _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_33 | _GEN_33; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_39 = _T_33 ? 2'h2 : _GEN_35; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_40 = _T_33 ? 2'h1 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_33 ? 1'h0 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_33 ? 1'h0 : _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_32 | _GEN_38; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_44 = _T_32 ? 2'h1 : _GEN_39; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_45 = _T_32 ? 2'h1 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_46 = _T_32 ? 1'h0 : _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_32 ? 1'h0 : _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_21 | _GEN_43; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_49 = _T_21 ? _GEN_26 : 4'h0; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_50 = _T_21 ? 2'h0 : _GEN_44; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_51 = _T_21 ? 2'h0 : _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_21 ? 1'h0 : _GEN_46; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_21 ? 1'h0 : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_11 | _GEN_48; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_55 = _T_11 ? 2'h1 : _GEN_51; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_56 = _T_11 ? _GEN_16 : _GEN_49; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_57 = _T_11 ? 2'h0 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_11 ? 1'h0 : _GEN_52; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_11 ? 1'h0 : _GEN_53; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_60 = _T_7 ? 2'h1 : _GEN_55; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_61 = _T_7 ? _GEN_7 : 4'h0; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_7 ? 1'h0 : _GEN_54; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_63 = _T_7 ? 4'h0 : _GEN_56; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_64 = _T_7 ? 2'h0 : _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_7 ? 1'h0 : _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_7 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_1 | _GEN_62; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_70 = _T_1 ? {{1'd0}, _GEN_4} : _GEN_61; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_71 = _T_1 ? 4'h0 : _GEN_63; // @[Conditional.scala 40:58]
  wire  _GEN_73 = _T_1 ? 1'h0 : _GEN_65; // @[Conditional.scala 40:58]
  RegFile regFile ( // @[ID.scala 21:23]
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_registerS1Index(regFile_io_registerS1Index),
    .io_registerS2Index(regFile_io_registerS2Index),
    .io_registerWIndex(regFile_io_registerWIndex),
    .io_registerWData(regFile_io_registerWData),
    .io_writeEn(regFile_io_writeEn),
    .io_registerS1Data(regFile_io_registerS1Data),
    .io_registerS2Data(regFile_io_registerS2Data)
  );
  ImmGen immGen ( // @[ID.scala 23:22]
    .io_instruction(immGen_io_instruction),
    .io_immediate(immGen_io_immediate)
  );
  assign out_pc = in_pc; // @[ID.scala 50:10]
  assign out_imm = immGen_io_immediate; // @[ID.scala 45:11]
  assign out_regOp1 = regFile_io_registerS1Data; // @[ID.scala 37:14]
  assign out_regOp2 = regFile_io_registerS2Data; // @[ID.scala 38:14]
  assign out_rs1 = in_instr[19:15]; // @[ID.scala 47:11]
  assign out_rs2 = in_instr[24:20]; // @[ID.scala 48:11]
  assign out_rd = in_instr[11:7]; // @[ID.scala 49:10]
  assign out_aluOp = ctrl_flushID ? 4'h0 : _GEN_71; // @[ID.scala 54:13 ID.scala 102:21 ID.scala 105:21 ID.scala 108:21 ID.scala 111:21 ID.scala 114:21 ID.scala 117:21 ID.scala 119:23 ID.scala 123:21 ID.scala 126:21 ID.scala 134:21 ID.scala 136:23 ID.scala 140:21 ID.scala 143:21 ID.scala 146:21 ID.scala 149:21 ID.scala 152:21 ID.scala 154:23 ID.scala 158:21 ID.scala 161:21 ID.scala 197:15]
  assign out_aluSrc1 = _T_1 ? 2'h0 : _GEN_64; // @[ID.scala 52:15 ID.scala 167:19 ID.scala 172:19 ID.scala 181:19 ID.scala 188:19]
  assign out_aluSrc2 = _T_1 ? 2'h1 : _GEN_60; // @[ID.scala 53:15 ID.scala 63:19 ID.scala 84:19 ID.scala 99:19 ID.scala 168:19 ID.scala 173:19 ID.scala 182:19 ID.scala 189:19]
  assign out_brSrc = _T_1 ? 1'h0 : _GEN_66; // @[ID.scala 58:13 ID.scala 187:17]
  assign out_pcSrc = ctrl_flushID ? 1'h0 : _GEN_73; // @[ID.scala 56:13 ID.scala 177:17 ID.scala 183:17 ID.scala 190:17 ID.scala 200:15]
  assign out_wb = ctrl_flushID ? 1'h0 : _GEN_67; // @[ID.scala 51:10 ID.scala 62:14 ID.scala 98:14 ID.scala 131:14 ID.scala 166:14 ID.scala 171:14 ID.scala 176:14 ID.scala 180:14 ID.scala 186:14 ID.scala 196:12]
  assign out_wbSrc = ctrl_flushID ? 1'h0 : _T_1; // @[ID.scala 57:13 ID.scala 64:17 ID.scala 199:15]
  assign out_mem = ctrl_flushID ? 4'h0 : _GEN_70; // @[ID.scala 55:11 ID.scala 67:19 ID.scala 70:19 ID.scala 73:19 ID.scala 76:19 ID.scala 79:19 ID.scala 87:19 ID.scala 90:19 ID.scala 93:19 ID.scala 198:13]
  assign out_jump = opcode[2]; // @[ID.scala 31:12]
  assign out_funct3 = in_instr[14:12]; // @[ID.scala 32:14]
  assign ctrl_instr = in_instr; // @[ID.scala 194:14]
  assign regFile_clock = clock;
  assign regFile_reset = reset;
  assign regFile_io_registerS1Index = in_instr[19:15]; // @[ID.scala 35:30]
  assign regFile_io_registerS2Index = in_instr[24:20]; // @[ID.scala 36:30]
  assign regFile_io_registerWIndex = wb_rd; // @[ID.scala 40:29]
  assign regFile_io_registerWData = wb_res; // @[ID.scala 41:28]
  assign regFile_io_writeEn = wb_wb; // @[ID.scala 42:22]
  assign immGen_io_instruction = in_instr; // @[ID.scala 44:25]
endmodule
module ALU(
  input  [31:0] io_source1,
  input  [31:0] io_source2,
  input  [3:0]  io_operation,
  output [31:0] io_output
);
  wire [31:0] _T_2 = $signed(io_source1) + $signed(io_source2); // @[ALU.scala 19:27]
  wire  _T_3 = 4'h1 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_6 = $signed(io_source1) - $signed(io_source2); // @[ALU.scala 23:31]
  wire  _T_7 = 4'h2 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_8 = io_source1; // @[ALU.scala 26:32]
  wire [62:0] _GEN_8 = {{31'd0}, _T_8}; // @[ALU.scala 26:39]
  wire [62:0] _T_11 = _GEN_8 << io_source2[4:0]; // @[ALU.scala 26:67]
  wire  _T_12 = 4'h3 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_16 = io_source1 >> io_source2[4:0]; // @[ALU.scala 29:67]
  wire  _T_17 = 4'h4 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_19 = $signed(io_source1) >>> io_source2[4:0]; // @[ALU.scala 32:32]
  wire  _T_20 = 4'h6 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_22 = $signed(io_source1) | $signed(io_source2); // @[ALU.scala 35:31]
  wire  _T_23 = 4'h5 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_25 = $signed(io_source1) & $signed(io_source2); // @[ALU.scala 38:31]
  wire  _T_26 = 4'h7 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_28 = $signed(io_source1) ^ $signed(io_source2); // @[ALU.scala 41:31]
  wire  _T_29 = 4'h8 == io_operation; // @[Conditional.scala 37:30]
  wire  _T_31 = $signed(io_source1) < $signed(io_source2); // @[ALU.scala 44:52]
  wire [31:0] _GEN_0 = _T_29 ? $signed({32{_T_31}}) : $signed(_T_2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1 = _T_26 ? $signed(_T_28) : $signed(_GEN_0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_23 ? $signed(_T_25) : $signed(_GEN_1); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_3 = _T_20 ? $signed(_T_22) : $signed(_GEN_2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_4 = _T_17 ? $signed(_T_19) : $signed(_GEN_3); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5 = _T_12 ? $signed(_T_16) : $signed(_GEN_4); // @[Conditional.scala 39:67]
  wire [62:0] _GEN_6 = _T_7 ? $signed(_T_11) : $signed({{31{_GEN_5[31]}},_GEN_5}); // @[Conditional.scala 39:67]
  wire [62:0] _GEN_7 = _T_3 ? $signed({{31{_T_6[31]}},_T_6}) : $signed(_GEN_6); // @[Conditional.scala 40:58]
  assign io_output = _GEN_7[31:0]; // @[ALU.scala 19:13 ALU.scala 23:17 ALU.scala 26:17 ALU.scala 29:17 ALU.scala 32:17 ALU.scala 35:17 ALU.scala 38:17 ALU.scala 41:17 ALU.scala 44:17]
endmodule
module BranchControl(
  input  [2:0]  io_funct3,
  input  [31:0] io_registerS1,
  input  [31:0] io_registerS2,
  input         io_jump,
  output        io_takeBranch
);
  wire  equal = $signed(io_registerS1) == $signed(io_registerS2); // @[BranchControl.scala 15:29]
  wire  lessThan = $signed(io_registerS1) < $signed(io_registerS2); // @[BranchControl.scala 16:32]
  wire  lessThanU = io_registerS1 < io_registerS2; // @[BranchControl.scala 17:42]
  wire  _T_2 = 3'h0 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_4 = ~equal; // @[BranchControl.scala 26:24]
  wire  _T_5 = 3'h4 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h5 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_7 = ~lessThan; // @[BranchControl.scala 32:24]
  wire  _T_8 = 3'h6 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h7 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_10 = ~lessThanU; // @[BranchControl.scala 38:24]
  wire  _GEN_0 = _T_9 & _T_10; // @[Conditional.scala 39:67]
  wire  _GEN_1 = _T_8 ? lessThanU : _GEN_0; // @[Conditional.scala 39:67]
  wire  _GEN_2 = _T_6 ? _T_7 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_5 ? lessThan : _GEN_2; // @[Conditional.scala 39:67]
  wire  _GEN_4 = _T_3 ? _T_4 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_2 ? equal : _GEN_4; // @[Conditional.scala 40:58]
  assign io_takeBranch = io_jump | _GEN_5; // @[BranchControl.scala 19:17 BranchControl.scala 23:21 BranchControl.scala 26:21 BranchControl.scala 29:21 BranchControl.scala 32:21 BranchControl.scala 35:21 BranchControl.scala 38:21 BranchControl.scala 42:19]
endmodule
module EX(
  input  [31:0] in_pc,
  input  [31:0] in_imm,
  input  [31:0] in_regOp1,
  input  [31:0] in_regOp2,
  input  [4:0]  in_rs1,
  input  [4:0]  in_rs2,
  input  [4:0]  in_rd,
  input  [3:0]  in_aluOp,
  input  [1:0]  in_aluSrc1,
  input  [1:0]  in_aluSrc2,
  input         in_brSrc,
  input         in_pcSrc,
  input         in_wb,
  input         in_wbSrc,
  input  [3:0]  in_mem,
  input         in_jump,
  input  [2:0]  in_funct3,
  output [31:0] out_aluRes,
  output [31:0] out_regOp2,
  output [4:0]  out_rd,
  output        out_wb,
  output        out_wbSrc,
  output [3:0]  out_mem,
  output [4:0]  ctrl_rs1,
  output [4:0]  ctrl_rs2,
  output [4:0]  ctrl_rd,
  input  [31:0] ctrl_fwdA,
  input  [31:0] ctrl_fwdB,
  input         ctrl_fwdA_en,
  input         ctrl_fwdB_en,
  output [31:0] ctrl_branchOut_pcNext,
  output        ctrl_branchOut_branch
);
  wire [31:0] alu_io_source1; // @[EX.scala 31:19]
  wire [31:0] alu_io_source2; // @[EX.scala 31:19]
  wire [3:0] alu_io_operation; // @[EX.scala 31:19]
  wire [31:0] alu_io_output; // @[EX.scala 31:19]
  wire [2:0] branchControl_io_funct3; // @[EX.scala 32:29]
  wire [31:0] branchControl_io_registerS1; // @[EX.scala 32:29]
  wire [31:0] branchControl_io_registerS2; // @[EX.scala 32:29]
  wire  branchControl_io_jump; // @[EX.scala 32:29]
  wire  branchControl_io_takeBranch; // @[EX.scala 32:29]
  wire [31:0] fwdRegOp1 = ctrl_fwdA_en ? $signed(ctrl_fwdA) : $signed(in_regOp1); // @[EX.scala 33:22]
  wire [31:0] fwdRegOp2 = ctrl_fwdB_en ? $signed(ctrl_fwdB) : $signed(in_regOp2); // @[EX.scala 34:22]
  wire  _T = branchControl_io_takeBranch; // @[EX.scala 41:58]
  wire [31:0] _T_5 = $signed(fwdRegOp1) + $signed(in_imm); // @[EX.scala 42:72]
  wire [31:0] _T_10 = $signed(in_pc) + $signed(in_imm); // @[EX.scala 42:112]
  wire  _T_19 = 2'h0 == in_aluSrc1; // @[Conditional.scala 37:30]
  wire  _T_20 = 2'h1 == in_aluSrc1; // @[Conditional.scala 37:30]
  wire  _T_22 = 2'h2 == in_aluSrc1; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_1 = _T_22 ? $signed(32'sh0) : $signed(fwdRegOp1); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_20 ? $signed(in_pc) : $signed(_GEN_1); // @[Conditional.scala 39:67]
  wire  _T_23 = 2'h0 == in_aluSrc2; // @[Conditional.scala 37:30]
  wire  _T_24 = 2'h1 == in_aluSrc2; // @[Conditional.scala 37:30]
  wire  _T_25 = 2'h2 == in_aluSrc2; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_4 = _T_25 ? $signed(32'sh4) : $signed(fwdRegOp2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5 = _T_24 ? $signed(in_imm) : $signed(_GEN_4); // @[Conditional.scala 39:67]
  ALU alu ( // @[EX.scala 31:19]
    .io_source1(alu_io_source1),
    .io_source2(alu_io_source2),
    .io_operation(alu_io_operation),
    .io_output(alu_io_output)
  );
  BranchControl branchControl ( // @[EX.scala 32:29]
    .io_funct3(branchControl_io_funct3),
    .io_registerS1(branchControl_io_registerS1),
    .io_registerS2(branchControl_io_registerS2),
    .io_jump(branchControl_io_jump),
    .io_takeBranch(branchControl_io_takeBranch)
  );
  assign out_aluRes = alu_io_output; // @[EX.scala 76:14]
  assign out_regOp2 = ctrl_fwdB_en ? $signed(ctrl_fwdB) : $signed(in_regOp2); // @[EX.scala 77:14]
  assign out_rd = in_rd; // @[EX.scala 24:10 EX.scala 29:10]
  assign out_wb = in_wb; // @[EX.scala 26:10]
  assign out_wbSrc = in_wbSrc; // @[EX.scala 28:13]
  assign out_mem = in_mem; // @[EX.scala 27:11]
  assign ctrl_rs1 = in_rs1; // @[EX.scala 22:12]
  assign ctrl_rs2 = in_rs2; // @[EX.scala 23:12]
  assign ctrl_rd = in_rd; // @[EX.scala 25:11]
  assign ctrl_branchOut_pcNext = in_brSrc ? _T_5 : _T_10; // @[EX.scala 42:25 EX.scala 46:27]
  assign ctrl_branchOut_branch = _T & in_pcSrc; // @[EX.scala 41:25]
  assign alu_io_source1 = _T_19 ? $signed(fwdRegOp1) : $signed(_GEN_2); // @[EX.scala 49:18 EX.scala 55:22 EX.scala 58:22 EX.scala 61:22]
  assign alu_io_source2 = _T_23 ? $signed(fwdRegOp2) : $signed(_GEN_5); // @[EX.scala 50:18 EX.scala 66:22 EX.scala 69:22 EX.scala 72:22]
  assign alu_io_operation = in_aluOp; // @[EX.scala 51:20]
  assign branchControl_io_funct3 = in_funct3; // @[EX.scala 36:27]
  assign branchControl_io_registerS1 = ctrl_fwdA_en ? $signed(ctrl_fwdA) : $signed(in_regOp1); // @[EX.scala 38:31]
  assign branchControl_io_registerS2 = ctrl_fwdB_en ? $signed(ctrl_fwdB) : $signed(in_regOp2); // @[EX.scala 39:31]
  assign branchControl_io_jump = in_jump; // @[EX.scala 37:25]
endmodule
module MEM(
  input         clock,
  input  [31:0] in_aluRes,
  input  [31:0] in_regOp2,
  input  [4:0]  in_rd,
  input         in_wb,
  input         in_wbSrc,
  input  [3:0]  in_mem,
  output [31:0] out_memRes,
  output [31:0] out_aluRes,
  output [4:0]  out_rd,
  output        out_wb,
  output        out_wbSrc,
  output [31:0] dataBus_addr,
  input  [7:0]  dataBus_rdData_0,
  input  [7:0]  dataBus_rdData_1,
  input  [7:0]  dataBus_rdData_2,
  input  [7:0]  dataBus_rdData_3,
  output [7:0]  dataBus_wrData_0,
  output [7:0]  dataBus_wrData_1,
  output [7:0]  dataBus_wrData_2,
  output [7:0]  dataBus_wrData_3,
  output        dataBus_we_0,
  output        dataBus_we_1,
  output        dataBus_we_2,
  output        dataBus_we_3,
  output        dataBus_w,
  output [4:0]  ctrl_rd,
  output [31:0] ctrl_aluRes
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _T_4 = 2'h1 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _T_6 = 2'h2 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _T_8 = 2'h3 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _GEN_4 = _T_6 | _T_8; // @[Conditional.scala 39:67]
  wire  _GEN_6 = _T_6 ? 1'h0 : _T_8; // @[Conditional.scala 39:67]
  wire  _GEN_8 = _T_4 | _GEN_4; // @[Conditional.scala 40:58]
  wire  _GEN_9 = _T_4 ? 1'h0 : _GEN_4; // @[Conditional.scala 40:58]
  wire  _GEN_10 = _T_4 ? 1'h0 : _GEN_6; // @[Conditional.scala 40:58]
  wire [31:0] _T_11 = in_regOp2; // @[MEM.scala 36:41]
  wire  _T_21 = in_mem[2] & dataBus_rdData_0[7]; // @[MEM.scala 43:56]
  wire [5:0] _T_96 = {_T_21,_T_21,_T_21,_T_21,_T_21,_T_21}; // @[MEM.scala 43:73]
  wire [11:0] _T_102 = {_T_21,_T_21,_T_21,_T_21,_T_21,_T_21,_T_96}; // @[MEM.scala 43:73]
  wire [31:0] _T_116 = {_T_21,_T_21,_T_21,_T_21,_T_21,_T_21,_T_96,_T_102,dataBus_rdData_0}; // @[MEM.scala 43:92]
  wire  _T_120 = in_mem[2] & dataBus_rdData_1[7]; // @[MEM.scala 46:56]
  wire [7:0] _T_173 = {_T_120,_T_120,_T_120,_T_120,_T_120,_T_120,_T_120,_T_120}; // @[MEM.scala 46:73]
  wire [23:0] _T_182 = {_T_120,_T_120,_T_120,_T_120,_T_120,_T_120,_T_120,_T_120,_T_173,dataBus_rdData_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_184 = {_T_182,dataBus_rdData_0}; // @[MEM.scala 46:103]
  wire [31:0] _T_189 = {dataBus_rdData_3,dataBus_rdData_2,dataBus_rdData_1,dataBus_rdData_0}; // @[MEM.scala 49:72]
  wire [31:0] _GEN_16 = _T_8 ? $signed(_T_189) : $signed(32'sh0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_17 = _T_6 ? $signed(_T_184) : $signed(_GEN_16); // @[Conditional.scala 39:67]
  reg [31:0] delayedAluRes; // @[MEM.scala 53:30]
  assign out_memRes = _T_4 ? $signed(_T_116) : $signed(_GEN_17); // @[MEM.scala 40:14 MEM.scala 43:18 MEM.scala 46:18 MEM.scala 49:18]
  assign out_aluRes = delayedAluRes; // @[MEM.scala 58:14]
  assign out_rd = in_rd; // @[MEM.scala 57:10]
  assign out_wb = in_wb; // @[MEM.scala 55:10]
  assign out_wbSrc = in_wbSrc; // @[MEM.scala 56:13]
  assign dataBus_addr = in_aluRes; // @[MEM.scala 35:16]
  assign dataBus_wrData_0 = _T_11[7:0]; // @[MEM.scala 36:18]
  assign dataBus_wrData_1 = _T_11[15:8]; // @[MEM.scala 36:18]
  assign dataBus_wrData_2 = _T_11[23:16]; // @[MEM.scala 36:18]
  assign dataBus_wrData_3 = _T_11[31:24]; // @[MEM.scala 36:18]
  assign dataBus_we_0 = in_mem[3] & _GEN_8; // @[MEM.scala 20:14 MEM.scala 25:20 MEM.scala 28:20 MEM.scala 31:20]
  assign dataBus_we_1 = in_mem[3] & _GEN_9; // @[MEM.scala 20:14 MEM.scala 25:20 MEM.scala 28:20 MEM.scala 31:20]
  assign dataBus_we_2 = in_mem[3] & _GEN_10; // @[MEM.scala 20:14 MEM.scala 25:20 MEM.scala 28:20 MEM.scala 31:20]
  assign dataBus_we_3 = in_mem[3] & _GEN_10; // @[MEM.scala 20:14 MEM.scala 25:20 MEM.scala 28:20 MEM.scala 31:20]
  assign dataBus_w = in_mem[3]; // @[MEM.scala 21:13]
  assign ctrl_rd = in_rd; // @[MEM.scala 60:11]
  assign ctrl_aluRes = delayedAluRes; // @[MEM.scala 59:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delayedAluRes = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    delayedAluRes <= in_aluRes;
  end
endmodule
module WB(
  input  [31:0] in_memRes,
  input  [31:0] in_aluRes,
  input  [4:0]  in_rd,
  input         in_wb,
  input         in_wbSrc,
  output [4:0]  out_rd,
  output [31:0] out_res,
  output        out_wb,
  output [4:0]  ctrl_rd,
  output [31:0] ctrl_res
);
  assign out_rd = in_rd; // @[WB.scala 17:10]
  assign out_res = in_wbSrc ? $signed(in_memRes) : $signed(in_aluRes); // @[WB.scala 14:11]
  assign out_wb = in_wb; // @[WB.scala 18:10]
  assign ctrl_rd = in_rd; // @[WB.scala 15:11]
  assign ctrl_res = in_wbSrc ? $signed(in_memRes) : $signed(in_aluRes); // @[WB.scala 16:12]
endmodule
module ForwardingUnit(
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd_MEM,
  input         io_wb_MEM,
  input  [4:0]  io_rd_WB,
  input         io_wb_WB,
  input  [31:0] io_aluRes_MEM,
  input  [31:0] io_res_WB,
  output [31:0] io_fwdA,
  output [31:0] io_fwdB,
  output        io_fwdA_en,
  output        io_fwdB_en
);
  wire  _T = io_rs1 == io_rd_MEM; // @[ForwardingUnit.scala 24:15]
  wire  _T_1 = _T & io_wb_MEM; // @[ForwardingUnit.scala 24:29]
  wire  _T_2 = io_rs1 == io_rd_WB; // @[ForwardingUnit.scala 28:21]
  wire  _T_3 = _T_2 & io_wb_WB; // @[ForwardingUnit.scala 28:34]
  wire [31:0] _GEN_1 = _T_3 ? $signed(io_res_WB) : $signed(32'sh0); // @[ForwardingUnit.scala 28:47]
  wire  _T_4 = io_rs2 == io_rd_MEM; // @[ForwardingUnit.scala 36:15]
  wire  _T_5 = _T_4 & io_wb_MEM; // @[ForwardingUnit.scala 36:29]
  wire  _T_6 = io_rs2 == io_rd_WB; // @[ForwardingUnit.scala 40:21]
  wire  _T_7 = _T_6 & io_wb_WB; // @[ForwardingUnit.scala 40:34]
  wire [31:0] _GEN_5 = _T_7 ? $signed(io_res_WB) : $signed(32'sh0); // @[ForwardingUnit.scala 40:47]
  assign io_fwdA = _T_1 ? $signed(io_aluRes_MEM) : $signed(_GEN_1); // @[ForwardingUnit.scala 26:13 ForwardingUnit.scala 30:13 ForwardingUnit.scala 32:13]
  assign io_fwdB = _T_5 ? $signed(io_aluRes_MEM) : $signed(_GEN_5); // @[ForwardingUnit.scala 38:13 ForwardingUnit.scala 42:13 ForwardingUnit.scala 44:13]
  assign io_fwdA_en = _T_1 | _T_3; // @[ForwardingUnit.scala 22:14 ForwardingUnit.scala 25:16 ForwardingUnit.scala 29:16]
  assign io_fwdB_en = _T_5 | _T_7; // @[ForwardingUnit.scala 35:14 ForwardingUnit.scala 37:16 ForwardingUnit.scala 41:16]
endmodule
module HazardDetectionUnit(
  output        io_pcEn,
  output        io_flushIF,
  output        io_flushID,
  output        io_enableIF_ID,
  input  [4:0]  io_rd_EX,
  input  [31:0] io_instr,
  input         io_wbSrc_EX,
  input         io_branch_EX
);
  wire [4:0] rs1 = io_instr[19:15]; // @[HazardDetectionUnit.scala 22:21]
  wire [4:0] rs2 = io_instr[24:20]; // @[HazardDetectionUnit.scala 23:21]
  wire  rs1IsAccessed = io_rd_EX == rs1; // @[HazardDetectionUnit.scala 24:32]
  wire  rs2IsAccessed = io_rd_EX == rs2; // @[HazardDetectionUnit.scala 25:32]
  wire  _T = rs1IsAccessed | rs2IsAccessed; // @[HazardDetectionUnit.scala 26:23]
  wire  _T_1 = _T & io_wbSrc_EX; // @[HazardDetectionUnit.scala 26:41]
  wire  _GEN_0 = _T_1 ? 1'h0 : 1'h1; // @[HazardDetectionUnit.scala 26:57]
  assign io_pcEn = _T_1 ? 1'h0 : 1'h1; // @[HazardDetectionUnit.scala 17:11 HazardDetectionUnit.scala 27:13]
  assign io_flushIF = io_branch_EX; // @[HazardDetectionUnit.scala 18:14 HazardDetectionUnit.scala 33:16]
  assign io_flushID = io_branch_EX | _T_1; // @[HazardDetectionUnit.scala 19:14 HazardDetectionUnit.scala 28:16 HazardDetectionUnit.scala 34:16]
  assign io_enableIF_ID = io_branch_EX ? 1'h0 : _GEN_0; // @[HazardDetectionUnit.scala 20:18 HazardDetectionUnit.scala 29:20 HazardDetectionUnit.scala 35:20]
endmodule
module RVCore(
  input         clock,
  input         reset,
  output [31:0] io_dataBus_addr,
  input  [7:0]  io_dataBus_rdData_0,
  input  [7:0]  io_dataBus_rdData_1,
  input  [7:0]  io_dataBus_rdData_2,
  input  [7:0]  io_dataBus_rdData_3,
  output [7:0]  io_dataBus_wrData_0,
  output [7:0]  io_dataBus_wrData_1,
  output [7:0]  io_dataBus_wrData_2,
  output [7:0]  io_dataBus_wrData_3,
  output        io_dataBus_we_0,
  output        io_dataBus_we_1,
  output        io_dataBus_we_2,
  output        io_dataBus_we_3,
  output        io_dataBus_w
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  ifStage_clock; // @[RVCore.scala 18:23]
  wire  ifStage_reset; // @[RVCore.scala 18:23]
  wire [31:0] ifStage_in_pcNext; // @[RVCore.scala 18:23]
  wire  ifStage_in_branch; // @[RVCore.scala 18:23]
  wire [31:0] ifStage_out_pc; // @[RVCore.scala 18:23]
  wire [31:0] ifStage_out_instr; // @[RVCore.scala 18:23]
  wire  ifStage_ctrl_pcEn; // @[RVCore.scala 18:23]
  wire  idStage_clock; // @[RVCore.scala 19:23]
  wire  idStage_reset; // @[RVCore.scala 19:23]
  wire [31:0] idStage_in_pc; // @[RVCore.scala 19:23]
  wire [31:0] idStage_in_instr; // @[RVCore.scala 19:23]
  wire [31:0] idStage_out_pc; // @[RVCore.scala 19:23]
  wire [31:0] idStage_out_imm; // @[RVCore.scala 19:23]
  wire [31:0] idStage_out_regOp1; // @[RVCore.scala 19:23]
  wire [31:0] idStage_out_regOp2; // @[RVCore.scala 19:23]
  wire [4:0] idStage_out_rs1; // @[RVCore.scala 19:23]
  wire [4:0] idStage_out_rs2; // @[RVCore.scala 19:23]
  wire [4:0] idStage_out_rd; // @[RVCore.scala 19:23]
  wire [3:0] idStage_out_aluOp; // @[RVCore.scala 19:23]
  wire [1:0] idStage_out_aluSrc1; // @[RVCore.scala 19:23]
  wire [1:0] idStage_out_aluSrc2; // @[RVCore.scala 19:23]
  wire  idStage_out_brSrc; // @[RVCore.scala 19:23]
  wire  idStage_out_pcSrc; // @[RVCore.scala 19:23]
  wire  idStage_out_wb; // @[RVCore.scala 19:23]
  wire  idStage_out_wbSrc; // @[RVCore.scala 19:23]
  wire [3:0] idStage_out_mem; // @[RVCore.scala 19:23]
  wire  idStage_out_jump; // @[RVCore.scala 19:23]
  wire [2:0] idStage_out_funct3; // @[RVCore.scala 19:23]
  wire [4:0] idStage_wb_rd; // @[RVCore.scala 19:23]
  wire [31:0] idStage_wb_res; // @[RVCore.scala 19:23]
  wire  idStage_wb_wb; // @[RVCore.scala 19:23]
  wire  idStage_ctrl_flushID; // @[RVCore.scala 19:23]
  wire [31:0] idStage_ctrl_instr; // @[RVCore.scala 19:23]
  wire [31:0] exStage_in_pc; // @[RVCore.scala 20:23]
  wire [31:0] exStage_in_imm; // @[RVCore.scala 20:23]
  wire [31:0] exStage_in_regOp1; // @[RVCore.scala 20:23]
  wire [31:0] exStage_in_regOp2; // @[RVCore.scala 20:23]
  wire [4:0] exStage_in_rs1; // @[RVCore.scala 20:23]
  wire [4:0] exStage_in_rs2; // @[RVCore.scala 20:23]
  wire [4:0] exStage_in_rd; // @[RVCore.scala 20:23]
  wire [3:0] exStage_in_aluOp; // @[RVCore.scala 20:23]
  wire [1:0] exStage_in_aluSrc1; // @[RVCore.scala 20:23]
  wire [1:0] exStage_in_aluSrc2; // @[RVCore.scala 20:23]
  wire  exStage_in_brSrc; // @[RVCore.scala 20:23]
  wire  exStage_in_pcSrc; // @[RVCore.scala 20:23]
  wire  exStage_in_wb; // @[RVCore.scala 20:23]
  wire  exStage_in_wbSrc; // @[RVCore.scala 20:23]
  wire [3:0] exStage_in_mem; // @[RVCore.scala 20:23]
  wire  exStage_in_jump; // @[RVCore.scala 20:23]
  wire [2:0] exStage_in_funct3; // @[RVCore.scala 20:23]
  wire [31:0] exStage_out_aluRes; // @[RVCore.scala 20:23]
  wire [31:0] exStage_out_regOp2; // @[RVCore.scala 20:23]
  wire [4:0] exStage_out_rd; // @[RVCore.scala 20:23]
  wire  exStage_out_wb; // @[RVCore.scala 20:23]
  wire  exStage_out_wbSrc; // @[RVCore.scala 20:23]
  wire [3:0] exStage_out_mem; // @[RVCore.scala 20:23]
  wire [4:0] exStage_ctrl_rs1; // @[RVCore.scala 20:23]
  wire [4:0] exStage_ctrl_rs2; // @[RVCore.scala 20:23]
  wire [4:0] exStage_ctrl_rd; // @[RVCore.scala 20:23]
  wire [31:0] exStage_ctrl_fwdA; // @[RVCore.scala 20:23]
  wire [31:0] exStage_ctrl_fwdB; // @[RVCore.scala 20:23]
  wire  exStage_ctrl_fwdA_en; // @[RVCore.scala 20:23]
  wire  exStage_ctrl_fwdB_en; // @[RVCore.scala 20:23]
  wire [31:0] exStage_ctrl_branchOut_pcNext; // @[RVCore.scala 20:23]
  wire  exStage_ctrl_branchOut_branch; // @[RVCore.scala 20:23]
  wire  memStage_clock; // @[RVCore.scala 21:24]
  wire [31:0] memStage_in_aluRes; // @[RVCore.scala 21:24]
  wire [31:0] memStage_in_regOp2; // @[RVCore.scala 21:24]
  wire [4:0] memStage_in_rd; // @[RVCore.scala 21:24]
  wire  memStage_in_wb; // @[RVCore.scala 21:24]
  wire  memStage_in_wbSrc; // @[RVCore.scala 21:24]
  wire [3:0] memStage_in_mem; // @[RVCore.scala 21:24]
  wire [31:0] memStage_out_memRes; // @[RVCore.scala 21:24]
  wire [31:0] memStage_out_aluRes; // @[RVCore.scala 21:24]
  wire [4:0] memStage_out_rd; // @[RVCore.scala 21:24]
  wire  memStage_out_wb; // @[RVCore.scala 21:24]
  wire  memStage_out_wbSrc; // @[RVCore.scala 21:24]
  wire [31:0] memStage_dataBus_addr; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_rdData_0; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_rdData_1; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_rdData_2; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_rdData_3; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_wrData_0; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_wrData_1; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_wrData_2; // @[RVCore.scala 21:24]
  wire [7:0] memStage_dataBus_wrData_3; // @[RVCore.scala 21:24]
  wire  memStage_dataBus_we_0; // @[RVCore.scala 21:24]
  wire  memStage_dataBus_we_1; // @[RVCore.scala 21:24]
  wire  memStage_dataBus_we_2; // @[RVCore.scala 21:24]
  wire  memStage_dataBus_we_3; // @[RVCore.scala 21:24]
  wire  memStage_dataBus_w; // @[RVCore.scala 21:24]
  wire [4:0] memStage_ctrl_rd; // @[RVCore.scala 21:24]
  wire [31:0] memStage_ctrl_aluRes; // @[RVCore.scala 21:24]
  wire [31:0] wbStage_in_memRes; // @[RVCore.scala 22:23]
  wire [31:0] wbStage_in_aluRes; // @[RVCore.scala 22:23]
  wire [4:0] wbStage_in_rd; // @[RVCore.scala 22:23]
  wire  wbStage_in_wb; // @[RVCore.scala 22:23]
  wire  wbStage_in_wbSrc; // @[RVCore.scala 22:23]
  wire [4:0] wbStage_out_rd; // @[RVCore.scala 22:23]
  wire [31:0] wbStage_out_res; // @[RVCore.scala 22:23]
  wire  wbStage_out_wb; // @[RVCore.scala 22:23]
  wire [4:0] wbStage_ctrl_rd; // @[RVCore.scala 22:23]
  wire [31:0] wbStage_ctrl_res; // @[RVCore.scala 22:23]
  wire [4:0] forwardingUnit_io_rs1; // @[RVCore.scala 29:30]
  wire [4:0] forwardingUnit_io_rs2; // @[RVCore.scala 29:30]
  wire [4:0] forwardingUnit_io_rd_MEM; // @[RVCore.scala 29:30]
  wire  forwardingUnit_io_wb_MEM; // @[RVCore.scala 29:30]
  wire [4:0] forwardingUnit_io_rd_WB; // @[RVCore.scala 29:30]
  wire  forwardingUnit_io_wb_WB; // @[RVCore.scala 29:30]
  wire [31:0] forwardingUnit_io_aluRes_MEM; // @[RVCore.scala 29:30]
  wire [31:0] forwardingUnit_io_res_WB; // @[RVCore.scala 29:30]
  wire [31:0] forwardingUnit_io_fwdA; // @[RVCore.scala 29:30]
  wire [31:0] forwardingUnit_io_fwdB; // @[RVCore.scala 29:30]
  wire  forwardingUnit_io_fwdA_en; // @[RVCore.scala 29:30]
  wire  forwardingUnit_io_fwdB_en; // @[RVCore.scala 29:30]
  wire  hazardDetectionUnit_io_pcEn; // @[RVCore.scala 30:35]
  wire  hazardDetectionUnit_io_flushIF; // @[RVCore.scala 30:35]
  wire  hazardDetectionUnit_io_flushID; // @[RVCore.scala 30:35]
  wire  hazardDetectionUnit_io_enableIF_ID; // @[RVCore.scala 30:35]
  wire [4:0] hazardDetectionUnit_io_rd_EX; // @[RVCore.scala 30:35]
  wire [31:0] hazardDetectionUnit_io_instr; // @[RVCore.scala 30:35]
  wire  hazardDetectionUnit_io_wbSrc_EX; // @[RVCore.scala 30:35]
  wire  hazardDetectionUnit_io_branch_EX; // @[RVCore.scala 30:35]
  reg [31:0] if_id_pc; // @[RVCore.scala 32:22]
  reg [31:0] if_id_instr; // @[RVCore.scala 32:22]
  reg [31:0] id_ex_pc; // @[RVCore.scala 33:22]
  reg [31:0] id_ex_imm; // @[RVCore.scala 33:22]
  reg [31:0] id_ex_regOp1; // @[RVCore.scala 33:22]
  reg [31:0] id_ex_regOp2; // @[RVCore.scala 33:22]
  reg [4:0] id_ex_rs1; // @[RVCore.scala 33:22]
  reg [4:0] id_ex_rs2; // @[RVCore.scala 33:22]
  reg [4:0] id_ex_rd; // @[RVCore.scala 33:22]
  reg [3:0] id_ex_aluOp; // @[RVCore.scala 33:22]
  reg [1:0] id_ex_aluSrc1; // @[RVCore.scala 33:22]
  reg [1:0] id_ex_aluSrc2; // @[RVCore.scala 33:22]
  reg  id_ex_brSrc; // @[RVCore.scala 33:22]
  reg  id_ex_pcSrc; // @[RVCore.scala 33:22]
  reg  id_ex_wb; // @[RVCore.scala 33:22]
  reg  id_ex_wbSrc; // @[RVCore.scala 33:22]
  reg [3:0] id_ex_mem; // @[RVCore.scala 33:22]
  reg  id_ex_jump; // @[RVCore.scala 33:22]
  reg [2:0] id_ex_funct3; // @[RVCore.scala 33:22]
  reg [31:0] ex_mem_regOp2; // @[RVCore.scala 34:23]
  reg [4:0] ex_mem_rd; // @[RVCore.scala 34:23]
  reg  ex_mem_wb; // @[RVCore.scala 34:23]
  reg  ex_mem_wbSrc; // @[RVCore.scala 34:23]
  reg [3:0] ex_mem_mem; // @[RVCore.scala 34:23]
  reg [31:0] mem_wb_memRes; // @[RVCore.scala 35:23]
  reg [31:0] mem_wb_aluRes; // @[RVCore.scala 35:23]
  reg [4:0] mem_wb_rd; // @[RVCore.scala 35:23]
  reg  mem_wb_wb; // @[RVCore.scala 35:23]
  reg  mem_wb_wbSrc; // @[RVCore.scala 35:23]
  IF ifStage ( // @[RVCore.scala 18:23]
    .clock(ifStage_clock),
    .reset(ifStage_reset),
    .in_pcNext(ifStage_in_pcNext),
    .in_branch(ifStage_in_branch),
    .out_pc(ifStage_out_pc),
    .out_instr(ifStage_out_instr),
    .ctrl_pcEn(ifStage_ctrl_pcEn)
  );
  ID idStage ( // @[RVCore.scala 19:23]
    .clock(idStage_clock),
    .reset(idStage_reset),
    .in_pc(idStage_in_pc),
    .in_instr(idStage_in_instr),
    .out_pc(idStage_out_pc),
    .out_imm(idStage_out_imm),
    .out_regOp1(idStage_out_regOp1),
    .out_regOp2(idStage_out_regOp2),
    .out_rs1(idStage_out_rs1),
    .out_rs2(idStage_out_rs2),
    .out_rd(idStage_out_rd),
    .out_aluOp(idStage_out_aluOp),
    .out_aluSrc1(idStage_out_aluSrc1),
    .out_aluSrc2(idStage_out_aluSrc2),
    .out_brSrc(idStage_out_brSrc),
    .out_pcSrc(idStage_out_pcSrc),
    .out_wb(idStage_out_wb),
    .out_wbSrc(idStage_out_wbSrc),
    .out_mem(idStage_out_mem),
    .out_jump(idStage_out_jump),
    .out_funct3(idStage_out_funct3),
    .wb_rd(idStage_wb_rd),
    .wb_res(idStage_wb_res),
    .wb_wb(idStage_wb_wb),
    .ctrl_flushID(idStage_ctrl_flushID),
    .ctrl_instr(idStage_ctrl_instr)
  );
  EX exStage ( // @[RVCore.scala 20:23]
    .in_pc(exStage_in_pc),
    .in_imm(exStage_in_imm),
    .in_regOp1(exStage_in_regOp1),
    .in_regOp2(exStage_in_regOp2),
    .in_rs1(exStage_in_rs1),
    .in_rs2(exStage_in_rs2),
    .in_rd(exStage_in_rd),
    .in_aluOp(exStage_in_aluOp),
    .in_aluSrc1(exStage_in_aluSrc1),
    .in_aluSrc2(exStage_in_aluSrc2),
    .in_brSrc(exStage_in_brSrc),
    .in_pcSrc(exStage_in_pcSrc),
    .in_wb(exStage_in_wb),
    .in_wbSrc(exStage_in_wbSrc),
    .in_mem(exStage_in_mem),
    .in_jump(exStage_in_jump),
    .in_funct3(exStage_in_funct3),
    .out_aluRes(exStage_out_aluRes),
    .out_regOp2(exStage_out_regOp2),
    .out_rd(exStage_out_rd),
    .out_wb(exStage_out_wb),
    .out_wbSrc(exStage_out_wbSrc),
    .out_mem(exStage_out_mem),
    .ctrl_rs1(exStage_ctrl_rs1),
    .ctrl_rs2(exStage_ctrl_rs2),
    .ctrl_rd(exStage_ctrl_rd),
    .ctrl_fwdA(exStage_ctrl_fwdA),
    .ctrl_fwdB(exStage_ctrl_fwdB),
    .ctrl_fwdA_en(exStage_ctrl_fwdA_en),
    .ctrl_fwdB_en(exStage_ctrl_fwdB_en),
    .ctrl_branchOut_pcNext(exStage_ctrl_branchOut_pcNext),
    .ctrl_branchOut_branch(exStage_ctrl_branchOut_branch)
  );
  MEM memStage ( // @[RVCore.scala 21:24]
    .clock(memStage_clock),
    .in_aluRes(memStage_in_aluRes),
    .in_regOp2(memStage_in_regOp2),
    .in_rd(memStage_in_rd),
    .in_wb(memStage_in_wb),
    .in_wbSrc(memStage_in_wbSrc),
    .in_mem(memStage_in_mem),
    .out_memRes(memStage_out_memRes),
    .out_aluRes(memStage_out_aluRes),
    .out_rd(memStage_out_rd),
    .out_wb(memStage_out_wb),
    .out_wbSrc(memStage_out_wbSrc),
    .dataBus_addr(memStage_dataBus_addr),
    .dataBus_rdData_0(memStage_dataBus_rdData_0),
    .dataBus_rdData_1(memStage_dataBus_rdData_1),
    .dataBus_rdData_2(memStage_dataBus_rdData_2),
    .dataBus_rdData_3(memStage_dataBus_rdData_3),
    .dataBus_wrData_0(memStage_dataBus_wrData_0),
    .dataBus_wrData_1(memStage_dataBus_wrData_1),
    .dataBus_wrData_2(memStage_dataBus_wrData_2),
    .dataBus_wrData_3(memStage_dataBus_wrData_3),
    .dataBus_we_0(memStage_dataBus_we_0),
    .dataBus_we_1(memStage_dataBus_we_1),
    .dataBus_we_2(memStage_dataBus_we_2),
    .dataBus_we_3(memStage_dataBus_we_3),
    .dataBus_w(memStage_dataBus_w),
    .ctrl_rd(memStage_ctrl_rd),
    .ctrl_aluRes(memStage_ctrl_aluRes)
  );
  WB wbStage ( // @[RVCore.scala 22:23]
    .in_memRes(wbStage_in_memRes),
    .in_aluRes(wbStage_in_aluRes),
    .in_rd(wbStage_in_rd),
    .in_wb(wbStage_in_wb),
    .in_wbSrc(wbStage_in_wbSrc),
    .out_rd(wbStage_out_rd),
    .out_res(wbStage_out_res),
    .out_wb(wbStage_out_wb),
    .ctrl_rd(wbStage_ctrl_rd),
    .ctrl_res(wbStage_ctrl_res)
  );
  ForwardingUnit forwardingUnit ( // @[RVCore.scala 29:30]
    .io_rs1(forwardingUnit_io_rs1),
    .io_rs2(forwardingUnit_io_rs2),
    .io_rd_MEM(forwardingUnit_io_rd_MEM),
    .io_wb_MEM(forwardingUnit_io_wb_MEM),
    .io_rd_WB(forwardingUnit_io_rd_WB),
    .io_wb_WB(forwardingUnit_io_wb_WB),
    .io_aluRes_MEM(forwardingUnit_io_aluRes_MEM),
    .io_res_WB(forwardingUnit_io_res_WB),
    .io_fwdA(forwardingUnit_io_fwdA),
    .io_fwdB(forwardingUnit_io_fwdB),
    .io_fwdA_en(forwardingUnit_io_fwdA_en),
    .io_fwdB_en(forwardingUnit_io_fwdB_en)
  );
  HazardDetectionUnit hazardDetectionUnit ( // @[RVCore.scala 30:35]
    .io_pcEn(hazardDetectionUnit_io_pcEn),
    .io_flushIF(hazardDetectionUnit_io_flushIF),
    .io_flushID(hazardDetectionUnit_io_flushID),
    .io_enableIF_ID(hazardDetectionUnit_io_enableIF_ID),
    .io_rd_EX(hazardDetectionUnit_io_rd_EX),
    .io_instr(hazardDetectionUnit_io_instr),
    .io_wbSrc_EX(hazardDetectionUnit_io_wbSrc_EX),
    .io_branch_EX(hazardDetectionUnit_io_branch_EX)
  );
  assign io_dataBus_addr = memStage_dataBus_addr; // @[RVCore.scala 80:14]
  assign io_dataBus_wrData_0 = memStage_dataBus_wrData_0; // @[RVCore.scala 80:14]
  assign io_dataBus_wrData_1 = memStage_dataBus_wrData_1; // @[RVCore.scala 80:14]
  assign io_dataBus_wrData_2 = memStage_dataBus_wrData_2; // @[RVCore.scala 80:14]
  assign io_dataBus_wrData_3 = memStage_dataBus_wrData_3; // @[RVCore.scala 80:14]
  assign io_dataBus_we_0 = memStage_dataBus_we_0; // @[RVCore.scala 80:14]
  assign io_dataBus_we_1 = memStage_dataBus_we_1; // @[RVCore.scala 80:14]
  assign io_dataBus_we_2 = memStage_dataBus_we_2; // @[RVCore.scala 80:14]
  assign io_dataBus_we_3 = memStage_dataBus_we_3; // @[RVCore.scala 80:14]
  assign io_dataBus_w = memStage_dataBus_w; // @[RVCore.scala 80:14]
  assign ifStage_clock = clock;
  assign ifStage_reset = reset;
  assign ifStage_in_pcNext = exStage_ctrl_branchOut_pcNext; // @[RVCore.scala 38:14]
  assign ifStage_in_branch = exStage_ctrl_branchOut_branch; // @[RVCore.scala 38:14]
  assign ifStage_ctrl_pcEn = hazardDetectionUnit_io_pcEn; // @[RVCore.scala 39:21]
  assign idStage_clock = clock;
  assign idStage_reset = reset;
  assign idStage_in_pc = if_id_pc; // @[RVCore.scala 48:14]
  assign idStage_in_instr = if_id_instr; // @[RVCore.scala 48:14]
  assign idStage_wb_rd = wbStage_out_rd; // @[RVCore.scala 47:14]
  assign idStage_wb_res = wbStage_out_res; // @[RVCore.scala 47:14]
  assign idStage_wb_wb = wbStage_out_wb; // @[RVCore.scala 47:14]
  assign idStage_ctrl_flushID = hazardDetectionUnit_io_flushID; // @[RVCore.scala 46:24]
  assign exStage_in_pc = id_ex_pc; // @[RVCore.scala 53:14]
  assign exStage_in_imm = id_ex_imm; // @[RVCore.scala 53:14]
  assign exStage_in_regOp1 = id_ex_regOp1; // @[RVCore.scala 53:14]
  assign exStage_in_regOp2 = id_ex_regOp2; // @[RVCore.scala 53:14]
  assign exStage_in_rs1 = id_ex_rs1; // @[RVCore.scala 53:14]
  assign exStage_in_rs2 = id_ex_rs2; // @[RVCore.scala 53:14]
  assign exStage_in_rd = id_ex_rd; // @[RVCore.scala 53:14]
  assign exStage_in_aluOp = id_ex_aluOp; // @[RVCore.scala 53:14]
  assign exStage_in_aluSrc1 = id_ex_aluSrc1; // @[RVCore.scala 53:14]
  assign exStage_in_aluSrc2 = id_ex_aluSrc2; // @[RVCore.scala 53:14]
  assign exStage_in_brSrc = id_ex_brSrc; // @[RVCore.scala 53:14]
  assign exStage_in_pcSrc = id_ex_pcSrc; // @[RVCore.scala 53:14]
  assign exStage_in_wb = id_ex_wb; // @[RVCore.scala 53:14]
  assign exStage_in_wbSrc = id_ex_wbSrc; // @[RVCore.scala 53:14]
  assign exStage_in_mem = id_ex_mem; // @[RVCore.scala 53:14]
  assign exStage_in_jump = id_ex_jump; // @[RVCore.scala 53:14]
  assign exStage_in_funct3 = id_ex_funct3; // @[RVCore.scala 53:14]
  assign exStage_ctrl_fwdA = forwardingUnit_io_fwdA; // @[RVCore.scala 60:21]
  assign exStage_ctrl_fwdB = forwardingUnit_io_fwdB; // @[RVCore.scala 61:21]
  assign exStage_ctrl_fwdA_en = forwardingUnit_io_fwdA_en; // @[RVCore.scala 62:24]
  assign exStage_ctrl_fwdB_en = forwardingUnit_io_fwdB_en; // @[RVCore.scala 63:24]
  assign memStage_clock = clock;
  assign memStage_in_aluRes = exStage_out_aluRes; // @[RVCore.scala 67:15 RVCore.scala 68:22]
  assign memStage_in_regOp2 = ex_mem_regOp2; // @[RVCore.scala 67:15]
  assign memStage_in_rd = ex_mem_rd; // @[RVCore.scala 67:15]
  assign memStage_in_wb = ex_mem_wb; // @[RVCore.scala 67:15]
  assign memStage_in_wbSrc = ex_mem_wbSrc; // @[RVCore.scala 67:15]
  assign memStage_in_mem = ex_mem_mem; // @[RVCore.scala 67:15]
  assign memStage_dataBus_rdData_0 = io_dataBus_rdData_0; // @[RVCore.scala 80:14]
  assign memStage_dataBus_rdData_1 = io_dataBus_rdData_1; // @[RVCore.scala 80:14]
  assign memStage_dataBus_rdData_2 = io_dataBus_rdData_2; // @[RVCore.scala 80:14]
  assign memStage_dataBus_rdData_3 = io_dataBus_rdData_3; // @[RVCore.scala 80:14]
  assign wbStage_in_memRes = mem_wb_memRes; // @[RVCore.scala 75:14]
  assign wbStage_in_aluRes = mem_wb_aluRes; // @[RVCore.scala 75:14]
  assign wbStage_in_rd = mem_wb_rd; // @[RVCore.scala 75:14]
  assign wbStage_in_wb = mem_wb_wb; // @[RVCore.scala 75:14]
  assign wbStage_in_wbSrc = mem_wb_wbSrc; // @[RVCore.scala 75:14]
  assign forwardingUnit_io_rs1 = exStage_ctrl_rs1; // @[RVCore.scala 55:25]
  assign forwardingUnit_io_rs2 = exStage_ctrl_rs2; // @[RVCore.scala 56:25]
  assign forwardingUnit_io_rd_MEM = memStage_ctrl_rd; // @[RVCore.scala 70:28]
  assign forwardingUnit_io_wb_MEM = memStage_out_wb; // @[RVCore.scala 72:28]
  assign forwardingUnit_io_rd_WB = wbStage_ctrl_rd; // @[RVCore.scala 76:27]
  assign forwardingUnit_io_wb_WB = wbStage_out_wb; // @[RVCore.scala 78:27]
  assign forwardingUnit_io_aluRes_MEM = memStage_ctrl_aluRes; // @[RVCore.scala 71:32]
  assign forwardingUnit_io_res_WB = wbStage_ctrl_res; // @[RVCore.scala 77:28]
  assign hazardDetectionUnit_io_rd_EX = exStage_ctrl_rd; // @[RVCore.scala 57:32]
  assign hazardDetectionUnit_io_instr = idStage_ctrl_instr; // @[RVCore.scala 45:32]
  assign hazardDetectionUnit_io_wbSrc_EX = exStage_out_wbSrc; // @[RVCore.scala 59:35]
  assign hazardDetectionUnit_io_branch_EX = exStage_ctrl_branchOut_branch; // @[RVCore.scala 58:36]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_id_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  if_id_instr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  id_ex_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  id_ex_imm = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  id_ex_regOp1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  id_ex_regOp2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  id_ex_rs1 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  id_ex_rs2 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  id_ex_rd = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  id_ex_aluOp = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  id_ex_aluSrc1 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  id_ex_aluSrc2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  id_ex_brSrc = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  id_ex_pcSrc = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  id_ex_wb = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  id_ex_wbSrc = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  id_ex_mem = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  id_ex_jump = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  id_ex_funct3 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  ex_mem_regOp2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  ex_mem_rd = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  ex_mem_wb = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ex_mem_wbSrc = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ex_mem_mem = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  mem_wb_memRes = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_wb_aluRes = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_wb_rd = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  mem_wb_wb = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mem_wb_wbSrc = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      if_id_pc <= 32'h0;
    end else if (hazardDetectionUnit_io_flushIF) begin
      if_id_pc <= 32'h0;
    end else if (hazardDetectionUnit_io_enableIF_ID) begin
      if_id_pc <= ifStage_out_pc;
    end
    if (reset) begin
      if_id_instr <= 32'sh0;
    end else if (hazardDetectionUnit_io_flushIF) begin
      if_id_instr <= 32'sh0;
    end else if (hazardDetectionUnit_io_enableIF_ID) begin
      if_id_instr <= ifStage_out_instr;
    end
    if (reset) begin
      id_ex_pc <= 32'h0;
    end else begin
      id_ex_pc <= idStage_out_pc;
    end
    if (reset) begin
      id_ex_imm <= 32'sh0;
    end else begin
      id_ex_imm <= idStage_out_imm;
    end
    if (reset) begin
      id_ex_regOp1 <= 32'sh0;
    end else begin
      id_ex_regOp1 <= idStage_out_regOp1;
    end
    if (reset) begin
      id_ex_regOp2 <= 32'sh0;
    end else begin
      id_ex_regOp2 <= idStage_out_regOp2;
    end
    if (reset) begin
      id_ex_rs1 <= 5'h0;
    end else begin
      id_ex_rs1 <= idStage_out_rs1;
    end
    if (reset) begin
      id_ex_rs2 <= 5'h0;
    end else begin
      id_ex_rs2 <= idStage_out_rs2;
    end
    if (reset) begin
      id_ex_rd <= 5'h0;
    end else begin
      id_ex_rd <= idStage_out_rd;
    end
    if (reset) begin
      id_ex_aluOp <= 4'h0;
    end else begin
      id_ex_aluOp <= idStage_out_aluOp;
    end
    if (reset) begin
      id_ex_aluSrc1 <= 2'h0;
    end else begin
      id_ex_aluSrc1 <= idStage_out_aluSrc1;
    end
    if (reset) begin
      id_ex_aluSrc2 <= 2'h0;
    end else begin
      id_ex_aluSrc2 <= idStage_out_aluSrc2;
    end
    if (reset) begin
      id_ex_brSrc <= 1'h0;
    end else begin
      id_ex_brSrc <= idStage_out_brSrc;
    end
    if (reset) begin
      id_ex_pcSrc <= 1'h0;
    end else begin
      id_ex_pcSrc <= idStage_out_pcSrc;
    end
    if (reset) begin
      id_ex_wb <= 1'h0;
    end else begin
      id_ex_wb <= idStage_out_wb;
    end
    if (reset) begin
      id_ex_wbSrc <= 1'h0;
    end else begin
      id_ex_wbSrc <= idStage_out_wbSrc;
    end
    if (reset) begin
      id_ex_mem <= 4'h0;
    end else begin
      id_ex_mem <= idStage_out_mem;
    end
    if (reset) begin
      id_ex_jump <= 1'h0;
    end else begin
      id_ex_jump <= idStage_out_jump;
    end
    if (reset) begin
      id_ex_funct3 <= 3'h0;
    end else begin
      id_ex_funct3 <= idStage_out_funct3;
    end
    if (reset) begin
      ex_mem_regOp2 <= 32'sh0;
    end else begin
      ex_mem_regOp2 <= exStage_out_regOp2;
    end
    if (reset) begin
      ex_mem_rd <= 5'h0;
    end else begin
      ex_mem_rd <= exStage_out_rd;
    end
    if (reset) begin
      ex_mem_wb <= 1'h0;
    end else begin
      ex_mem_wb <= exStage_out_wb;
    end
    if (reset) begin
      ex_mem_wbSrc <= 1'h0;
    end else begin
      ex_mem_wbSrc <= exStage_out_wbSrc;
    end
    if (reset) begin
      ex_mem_mem <= 4'h0;
    end else begin
      ex_mem_mem <= exStage_out_mem;
    end
    if (reset) begin
      mem_wb_memRes <= 32'sh0;
    end else begin
      mem_wb_memRes <= memStage_out_memRes;
    end
    if (reset) begin
      mem_wb_aluRes <= 32'sh0;
    end else begin
      mem_wb_aluRes <= memStage_out_aluRes;
    end
    if (reset) begin
      mem_wb_rd <= 5'h0;
    end else begin
      mem_wb_rd <= memStage_out_rd;
    end
    if (reset) begin
      mem_wb_wb <= 1'h0;
    end else begin
      mem_wb_wb <= memStage_out_wb;
    end
    if (reset) begin
      mem_wb_wbSrc <= 1'h0;
    end else begin
      mem_wb_wbSrc <= memStage_out_wbSrc;
    end
  end
endmodule
module RingBuffer(
  input        clock,
  input        reset,
  input        io_enq_write,
  output       io_enq_full,
  input  [7:0] io_enq_data,
  input        io_deq_read,
  output       io_deq_empty,
  output [7:0] io_deq_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem_0; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_1; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_2; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_3; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_4; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_5; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_6; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_7; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_8; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_9; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_10; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_11; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_12; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_13; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_14; // @[RingBuffer.scala 14:20]
  reg [7:0] mem_15; // @[RingBuffer.scala 14:20]
  reg [3:0] head; // @[RingBuffer.scala 15:21]
  reg [3:0] tail; // @[RingBuffer.scala 16:21]
  reg  wrapBitHead; // @[RingBuffer.scala 17:28]
  reg  wrapBitTail; // @[RingBuffer.scala 18:28]
  wire  _T_1 = head == tail; // @[RingBuffer.scala 27:13]
  wire  _T_2 = wrapBitHead == wrapBitTail; // @[RingBuffer.scala 28:22]
  wire  _GEN_1 = _T_2 ? 1'h0 : 1'h1; // @[RingBuffer.scala 28:39]
  wire  empty = _T_1 & _T_2; // @[RingBuffer.scala 27:23]
  wire  full = _T_1 & _GEN_1; // @[RingBuffer.scala 27:23]
  wire  _T_3 = ~full; // @[RingBuffer.scala 36:24]
  wire  _T_4 = io_enq_write & _T_3; // @[RingBuffer.scala 36:21]
  wire  _T_5 = head == 4'hf; // @[RingBuffer.scala 38:15]
  wire  _T_6 = ~wrapBitHead; // @[RingBuffer.scala 40:22]
  wire [3:0] _T_8 = head + 4'h1; // @[RingBuffer.scala 42:20]
  wire [7:0] _GEN_41 = 4'h1 == tail ? mem_1 : mem_0; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_42 = 4'h2 == tail ? mem_2 : _GEN_41; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_43 = 4'h3 == tail ? mem_3 : _GEN_42; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_44 = 4'h4 == tail ? mem_4 : _GEN_43; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_45 = 4'h5 == tail ? mem_5 : _GEN_44; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_46 = 4'h6 == tail ? mem_6 : _GEN_45; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_47 = 4'h7 == tail ? mem_7 : _GEN_46; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_48 = 4'h8 == tail ? mem_8 : _GEN_47; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_49 = 4'h9 == tail ? mem_9 : _GEN_48; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_50 = 4'ha == tail ? mem_10 : _GEN_49; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_51 = 4'hb == tail ? mem_11 : _GEN_50; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_52 = 4'hc == tail ? mem_12 : _GEN_51; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_53 = 4'hd == tail ? mem_13 : _GEN_52; // @[RingBuffer.scala 47:15]
  wire [7:0] _GEN_54 = 4'he == tail ? mem_14 : _GEN_53; // @[RingBuffer.scala 47:15]
  wire  _T_9 = ~empty; // @[RingBuffer.scala 48:23]
  wire  _T_10 = io_deq_read & _T_9; // @[RingBuffer.scala 48:20]
  wire  _T_11 = tail == 4'hf; // @[RingBuffer.scala 49:15]
  wire  _T_12 = ~wrapBitTail; // @[RingBuffer.scala 51:22]
  wire [3:0] _T_14 = tail + 4'h1; // @[RingBuffer.scala 53:20]
  assign io_enq_full = _T_1 & _GEN_1; // @[RingBuffer.scala 57:15]
  assign io_deq_empty = _T_1 & _T_2; // @[RingBuffer.scala 58:16]
  assign io_deq_data = 4'hf == tail ? mem_15 : _GEN_54; // @[RingBuffer.scala 47:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  head = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  tail = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  wrapBitHead = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  wrapBitTail = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mem_0 <= 8'h0;
    end else if (_T_4) begin
      if (4'h0 == head) begin
        mem_0 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_1 <= 8'h0;
    end else if (_T_4) begin
      if (4'h1 == head) begin
        mem_1 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_2 <= 8'h0;
    end else if (_T_4) begin
      if (4'h2 == head) begin
        mem_2 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_3 <= 8'h0;
    end else if (_T_4) begin
      if (4'h3 == head) begin
        mem_3 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_4 <= 8'h0;
    end else if (_T_4) begin
      if (4'h4 == head) begin
        mem_4 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_5 <= 8'h0;
    end else if (_T_4) begin
      if (4'h5 == head) begin
        mem_5 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_6 <= 8'h0;
    end else if (_T_4) begin
      if (4'h6 == head) begin
        mem_6 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_7 <= 8'h0;
    end else if (_T_4) begin
      if (4'h7 == head) begin
        mem_7 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_8 <= 8'h0;
    end else if (_T_4) begin
      if (4'h8 == head) begin
        mem_8 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_9 <= 8'h0;
    end else if (_T_4) begin
      if (4'h9 == head) begin
        mem_9 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_10 <= 8'h0;
    end else if (_T_4) begin
      if (4'ha == head) begin
        mem_10 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_11 <= 8'h0;
    end else if (_T_4) begin
      if (4'hb == head) begin
        mem_11 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_12 <= 8'h0;
    end else if (_T_4) begin
      if (4'hc == head) begin
        mem_12 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_13 <= 8'h0;
    end else if (_T_4) begin
      if (4'hd == head) begin
        mem_13 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_14 <= 8'h0;
    end else if (_T_4) begin
      if (4'he == head) begin
        mem_14 <= io_enq_data;
      end
    end
    if (reset) begin
      mem_15 <= 8'h0;
    end else if (_T_4) begin
      if (4'hf == head) begin
        mem_15 <= io_enq_data;
      end
    end
    if (reset) begin
      head <= 4'h0;
    end else if (_T_4) begin
      if (_T_5) begin
        head <= 4'h0;
      end else begin
        head <= _T_8;
      end
    end
    if (reset) begin
      tail <= 4'h0;
    end else if (_T_10) begin
      if (_T_11) begin
        tail <= 4'h0;
      end else begin
        tail <= _T_14;
      end
    end
    if (reset) begin
      wrapBitHead <= 1'h0;
    end else if (_T_4) begin
      if (_T_5) begin
        wrapBitHead <= _T_6;
      end
    end
    if (reset) begin
      wrapBitTail <= 1'h0;
    end else if (_T_10) begin
      if (_T_11) begin
        wrapBitTail <= _T_12;
      end
    end
  end
endmodule
module PS2(
  input        clock,
  input        reset,
  input        ps2_clk,
  input        ps2_data,
  output [7:0] bus_data,
  output [7:0] bus_flag,
  input        bus_clear
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  buffer_clock; // @[PS2.scala 18:22]
  wire  buffer_reset; // @[PS2.scala 18:22]
  wire  buffer_io_enq_write; // @[PS2.scala 18:22]
  wire  buffer_io_enq_full; // @[PS2.scala 18:22]
  wire [7:0] buffer_io_enq_data; // @[PS2.scala 18:22]
  wire  buffer_io_deq_read; // @[PS2.scala 18:22]
  wire  buffer_io_deq_empty; // @[PS2.scala 18:22]
  wire [7:0] buffer_io_deq_data; // @[PS2.scala 18:22]
  reg [10:0] shiftReg; // @[PS2.scala 21:25]
  reg [3:0] countReg; // @[PS2.scala 22:25]
  wire [10:0] _T_1 = {ps2_data,shiftReg[10:1]}; // @[Cat.scala 29:58]
  wire  _T_3 = ~buffer_io_deq_empty; // @[PS2.scala 27:16]
  wire  _T_4 = ~ps2_clk; // @[PS2.scala 30:8]
  reg  _T_5; // @[PS2.scala 30:35]
  reg  _T_6; // @[PS2.scala 30:27]
  wire  _T_7 = _T_4 & _T_6; // @[PS2.scala 30:17]
  wire [3:0] _T_9 = countReg + 4'h1; // @[PS2.scala 31:26]
  wire  _T_12 = countReg >= 4'h9; // @[PS2.scala 33:19]
  wire  _T_13 = ~buffer_io_enq_full; // @[PS2.scala 35:12]
  wire  _GEN_2 = _T_12 & _T_13; // @[PS2.scala 33:26]
  RingBuffer buffer ( // @[PS2.scala 18:22]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .io_enq_write(buffer_io_enq_write),
    .io_enq_full(buffer_io_enq_full),
    .io_enq_data(buffer_io_enq_data),
    .io_deq_read(buffer_io_deq_read),
    .io_deq_empty(buffer_io_deq_empty),
    .io_deq_data(buffer_io_deq_data)
  );
  assign bus_data = buffer_io_deq_data; // @[PS2.scala 26:12]
  assign bus_flag = {{7'd0}, _T_3}; // @[PS2.scala 27:12]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_io_enq_write = _T_7 & _GEN_2; // @[PS2.scala 19:23 PS2.scala 36:29]
  assign buffer_io_enq_data = _T_1[8:1]; // @[PS2.scala 24:22]
  assign buffer_io_deq_read = bus_clear; // @[PS2.scala 28:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftReg = _RAND_0[10:0];
  _RAND_1 = {1{`RANDOM}};
  countReg = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _T_5 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_6 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      shiftReg <= 11'h0;
    end else if (_T_7) begin
      shiftReg <= _T_1;
    end
    if (reset) begin
      countReg <= 4'h0;
    end else if (_T_7) begin
      if (_T_12) begin
        countReg <= 4'h0;
      end else begin
        countReg <= _T_9;
      end
    end
    _T_5 <= ps2_clk;
    _T_6 <= _T_5;
  end
endmodule
module RAM(
  input         clock,
  input  [31:0] io_addr,
  output [7:0]  io_rdData_0,
  output [7:0]  io_rdData_1,
  output [7:0]  io_rdData_2,
  output [7:0]  io_rdData_3,
  input  [7:0]  io_wrData_0,
  input  [7:0]  io_wrData_1,
  input  [7:0]  io_wrData_2,
  input  [7:0]  io_wrData_3,
  input         io_we_0,
  input         io_we_1,
  input         io_we_2,
  input         io_we_3,
  input         io_w
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] banks_0 [0:1023]; // @[RAM.scala 9:30]
  wire [7:0] banks_0__T_9_data; // @[RAM.scala 9:30]
  wire [9:0] banks_0__T_9_addr; // @[RAM.scala 9:30]
  wire [7:0] banks_0__T_78_data; // @[RAM.scala 9:30]
  wire [9:0] banks_0__T_78_addr; // @[RAM.scala 9:30]
  wire  banks_0__T_78_mask; // @[RAM.scala 9:30]
  wire  banks_0__T_78_en; // @[RAM.scala 9:30]
  reg [7:0] banks_1 [0:1023]; // @[RAM.scala 9:30]
  wire [7:0] banks_1__T_18_data; // @[RAM.scala 9:30]
  wire [9:0] banks_1__T_18_addr; // @[RAM.scala 9:30]
  wire [7:0] banks_1__T_87_data; // @[RAM.scala 9:30]
  wire [9:0] banks_1__T_87_addr; // @[RAM.scala 9:30]
  wire  banks_1__T_87_mask; // @[RAM.scala 9:30]
  wire  banks_1__T_87_en; // @[RAM.scala 9:30]
  reg [7:0] banks_2 [0:1023]; // @[RAM.scala 9:30]
  wire [7:0] banks_2__T_27_data; // @[RAM.scala 9:30]
  wire [9:0] banks_2__T_27_addr; // @[RAM.scala 9:30]
  wire [7:0] banks_2__T_96_data; // @[RAM.scala 9:30]
  wire [9:0] banks_2__T_96_addr; // @[RAM.scala 9:30]
  wire  banks_2__T_96_mask; // @[RAM.scala 9:30]
  wire  banks_2__T_96_en; // @[RAM.scala 9:30]
  reg [7:0] banks_3 [0:1023]; // @[RAM.scala 9:30]
  wire [7:0] banks_3__T_36_data; // @[RAM.scala 9:30]
  wire [9:0] banks_3__T_36_addr; // @[RAM.scala 9:30]
  wire [7:0] banks_3__T_105_data; // @[RAM.scala 9:30]
  wire [9:0] banks_3__T_105_addr; // @[RAM.scala 9:30]
  wire  banks_3__T_105_mask; // @[RAM.scala 9:30]
  wire  banks_3__T_105_en; // @[RAM.scala 9:30]
  reg [31:0] address; // @[RAM.scala 11:24]
  wire [1:0] byteOffset = address[1:0]; // @[RAM.scala 14:24]
  wire  _T_2 = byteOffset > 2'h0; // @[RAM.scala 16:78]
  wire [29:0] _T_5 = address[31:2] + 30'h1; // @[RAM.scala 16:100]
  wire [29:0] _T_7 = _T_2 ? _T_5 : address[31:2]; // @[RAM.scala 16:63]
  wire  _T_11 = byteOffset > 2'h1; // @[RAM.scala 16:78]
  wire [29:0] _T_16 = _T_11 ? _T_5 : address[31:2]; // @[RAM.scala 16:63]
  wire  _T_20 = byteOffset > 2'h2; // @[RAM.scala 16:78]
  wire [29:0] _T_25 = _T_20 ? _T_5 : address[31:2]; // @[RAM.scala 16:63]
  wire [2:0] _T_37 = {{1'd0}, byteOffset}; // @[RAM.scala 17:64]
  wire [1:0] _T_40 = byteOffset + 2'h1; // @[RAM.scala 17:64]
  wire [1:0] _T_42 = byteOffset + 2'h2; // @[RAM.scala 17:64]
  wire [1:0] _T_44 = byteOffset + 2'h3; // @[RAM.scala 17:64]
  wire [7:0] rdPorts_0 = banks_0__T_9_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] rdPorts_1 = banks_1__T_18_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] _GEN_1 = 2'h1 == _T_37[1:0] ? rdPorts_1 : rdPorts_0; // @[RAM.scala 17:23]
  wire [7:0] rdPorts_2 = banks_2__T_27_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] _GEN_2 = 2'h2 == _T_37[1:0] ? rdPorts_2 : _GEN_1; // @[RAM.scala 17:23]
  wire [7:0] rdPorts_3 = banks_3__T_36_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] _GEN_5 = 2'h1 == _T_40 ? rdPorts_1 : rdPorts_0; // @[RAM.scala 17:23]
  wire [7:0] _GEN_6 = 2'h2 == _T_40 ? rdPorts_2 : _GEN_5; // @[RAM.scala 17:23]
  wire [7:0] _GEN_9 = 2'h1 == _T_42 ? rdPorts_1 : rdPorts_0; // @[RAM.scala 17:23]
  wire [7:0] _GEN_10 = 2'h2 == _T_42 ? rdPorts_2 : _GEN_9; // @[RAM.scala 17:23]
  wire [7:0] _GEN_13 = 2'h1 == _T_44 ? rdPorts_1 : rdPorts_0; // @[RAM.scala 17:23]
  wire [7:0] _GEN_14 = 2'h2 == _T_44 ? rdPorts_2 : _GEN_13; // @[RAM.scala 17:23]
  wire [31:0] wrData = {io_wrData_3,io_wrData_2,io_wrData_1,io_wrData_0}; // @[Cat.scala 29:58]
  wire [7:0] wrDataInVec_3 = wrData[7:0]; // @[RAM.scala 28:68]
  wire [7:0] wrDataInVec_2 = wrData[15:8]; // @[RAM.scala 28:68]
  wire [7:0] wrDataInVec_1 = wrData[23:16]; // @[RAM.scala 28:68]
  wire [7:0] wrDataInVec_0 = wrData[31:24]; // @[RAM.scala 28:68]
  wire [7:0] _GEN_17 = 2'h1 == _T_44 ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 29:34]
  wire [7:0] _GEN_18 = 2'h2 == _T_44 ? wrDataInVec_2 : _GEN_17; // @[RAM.scala 29:34]
  wire [7:0] _GEN_21 = 2'h1 == _T_42 ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 29:34]
  wire [7:0] _GEN_22 = 2'h2 == _T_42 ? wrDataInVec_2 : _GEN_21; // @[RAM.scala 29:34]
  wire [7:0] _GEN_25 = 2'h1 == _T_40 ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 29:34]
  wire [7:0] _GEN_26 = 2'h2 == _T_40 ? wrDataInVec_2 : _GEN_25; // @[RAM.scala 29:34]
  wire [7:0] _GEN_29 = 2'h1 == _T_37[1:0] ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 29:34]
  wire [7:0] _GEN_30 = 2'h2 == _T_37[1:0] ? wrDataInVec_2 : _GEN_29; // @[RAM.scala 29:34]
  wire  _GEN_33 = 2'h1 == _T_37[1:0] ? io_we_1 : io_we_0; // @[RAM.scala 30:22]
  wire  _GEN_34 = 2'h2 == _T_37[1:0] ? io_we_2 : _GEN_33; // @[RAM.scala 30:22]
  wire  enVec_0 = 2'h3 == _T_37[1:0] ? io_we_3 : _GEN_34; // @[RAM.scala 30:22]
  wire  _GEN_37 = 2'h1 == _T_40 ? io_we_1 : io_we_0; // @[RAM.scala 30:22]
  wire  _GEN_38 = 2'h2 == _T_40 ? io_we_2 : _GEN_37; // @[RAM.scala 30:22]
  wire  enVec_1 = 2'h3 == _T_40 ? io_we_3 : _GEN_38; // @[RAM.scala 30:22]
  wire  _GEN_41 = 2'h1 == _T_42 ? io_we_1 : io_we_0; // @[RAM.scala 30:22]
  wire  _GEN_42 = 2'h2 == _T_42 ? io_we_2 : _GEN_41; // @[RAM.scala 30:22]
  wire  enVec_2 = 2'h3 == _T_42 ? io_we_3 : _GEN_42; // @[RAM.scala 30:22]
  wire  _GEN_45 = 2'h1 == _T_44 ? io_we_1 : io_we_0; // @[RAM.scala 30:22]
  wire  _GEN_46 = 2'h2 == _T_44 ? io_we_2 : _GEN_45; // @[RAM.scala 30:22]
  wire  enVec_3 = 2'h3 == _T_44 ? io_we_3 : _GEN_46; // @[RAM.scala 30:22]
  assign banks_0__T_9_addr = _T_7[9:0];
  assign banks_0__T_9_data = banks_0[banks_0__T_9_addr]; // @[RAM.scala 9:30]
  assign banks_0__T_78_data = 2'h3 == _T_44 ? wrDataInVec_3 : _GEN_18;
  assign banks_0__T_78_addr = _T_7[9:0];
  assign banks_0__T_78_mask = 1'h1;
  assign banks_0__T_78_en = io_w & enVec_0;
  assign banks_1__T_18_addr = _T_16[9:0];
  assign banks_1__T_18_data = banks_1[banks_1__T_18_addr]; // @[RAM.scala 9:30]
  assign banks_1__T_87_data = 2'h3 == _T_42 ? wrDataInVec_3 : _GEN_22;
  assign banks_1__T_87_addr = _T_16[9:0];
  assign banks_1__T_87_mask = 1'h1;
  assign banks_1__T_87_en = io_w & enVec_1;
  assign banks_2__T_27_addr = _T_25[9:0];
  assign banks_2__T_27_data = banks_2[banks_2__T_27_addr]; // @[RAM.scala 9:30]
  assign banks_2__T_96_data = 2'h3 == _T_40 ? wrDataInVec_3 : _GEN_26;
  assign banks_2__T_96_addr = _T_25[9:0];
  assign banks_2__T_96_mask = 1'h1;
  assign banks_2__T_96_en = io_w & enVec_2;
  assign banks_3__T_36_addr = address[11:2];
  assign banks_3__T_36_data = banks_3[banks_3__T_36_addr]; // @[RAM.scala 9:30]
  assign banks_3__T_105_data = 2'h3 == _T_37[1:0] ? wrDataInVec_3 : _GEN_30;
  assign banks_3__T_105_addr = address[11:2];
  assign banks_3__T_105_mask = 1'h1;
  assign banks_3__T_105_en = io_w & enVec_3;
  assign io_rdData_0 = 2'h3 == _T_37[1:0] ? rdPorts_3 : _GEN_2; // @[RAM.scala 17:13]
  assign io_rdData_1 = 2'h3 == _T_40 ? rdPorts_3 : _GEN_6; // @[RAM.scala 17:13]
  assign io_rdData_2 = 2'h3 == _T_42 ? rdPorts_3 : _GEN_10; // @[RAM.scala 17:13]
  assign io_rdData_3 = 2'h3 == _T_44 ? rdPorts_3 : _GEN_14; // @[RAM.scala 17:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_0[initvar] = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_1[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_2[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_3[initvar] = _RAND_3[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  address = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(banks_0__T_78_en & banks_0__T_78_mask) begin
      banks_0[banks_0__T_78_addr] <= banks_0__T_78_data; // @[RAM.scala 9:30]
    end
    if(banks_1__T_87_en & banks_1__T_87_mask) begin
      banks_1[banks_1__T_87_addr] <= banks_1__T_87_data; // @[RAM.scala 9:30]
    end
    if(banks_2__T_96_en & banks_2__T_96_mask) begin
      banks_2[banks_2__T_96_addr] <= banks_2__T_96_data; // @[RAM.scala 9:30]
    end
    if(banks_3__T_105_en & banks_3__T_105_mask) begin
      banks_3[banks_3__T_105_addr] <= banks_3__T_105_data; // @[RAM.scala 9:30]
    end
    address <= io_addr;
  end
endmodule
module SevenSeg(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [3:0]  io_out_anode,
  output [6:0]  io_out_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] _T; // @[SevenSeg.scala 20:25]
  wire  ticker = _T == 19'h7a120; // @[SevenSeg.scala 21:23]
  wire [18:0] _T_2 = _T + 19'h1; // @[SevenSeg.scala 22:37]
  reg [1:0] sevAnCounter; // @[SevenSeg.scala 13:25]
  wire  _T_4 = sevAnCounter == 2'h3; // @[SevenSeg.scala 15:28]
  wire [1:0] _T_6 = sevAnCounter + 2'h1; // @[SevenSeg.scala 15:51]
  wire  _T_8 = 2'h0 == sevAnCounter; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_2 = 4'h1 == io_in[15:12] ? 7'h79 : 7'h40; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_3 = 4'h2 == io_in[15:12] ? 7'h24 : _GEN_2; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_4 = 4'h3 == io_in[15:12] ? 7'h30 : _GEN_3; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_5 = 4'h4 == io_in[15:12] ? 7'h19 : _GEN_4; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_6 = 4'h5 == io_in[15:12] ? 7'h12 : _GEN_5; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_7 = 4'h6 == io_in[15:12] ? 7'h2 : _GEN_6; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_8 = 4'h7 == io_in[15:12] ? 7'h78 : _GEN_7; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_9 = 4'h8 == io_in[15:12] ? 7'h0 : _GEN_8; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_10 = 4'h9 == io_in[15:12] ? 7'h10 : _GEN_9; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_11 = 4'ha == io_in[15:12] ? 7'h8 : _GEN_10; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_12 = 4'hb == io_in[15:12] ? 7'h3 : _GEN_11; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_13 = 4'hc == io_in[15:12] ? 7'h46 : _GEN_12; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_14 = 4'hd == io_in[15:12] ? 7'h21 : _GEN_13; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_15 = 4'he == io_in[15:12] ? 7'h6 : _GEN_14; // @[SevenSeg.scala 54:20]
  wire [6:0] _GEN_16 = 4'hf == io_in[15:12] ? 7'he : _GEN_15; // @[SevenSeg.scala 54:20]
  wire  _T_10 = 2'h1 == sevAnCounter; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_18 = 4'h1 == io_in[11:8] ? 7'h79 : 7'h40; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_19 = 4'h2 == io_in[11:8] ? 7'h24 : _GEN_18; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_20 = 4'h3 == io_in[11:8] ? 7'h30 : _GEN_19; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_21 = 4'h4 == io_in[11:8] ? 7'h19 : _GEN_20; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_22 = 4'h5 == io_in[11:8] ? 7'h12 : _GEN_21; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_23 = 4'h6 == io_in[11:8] ? 7'h2 : _GEN_22; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_24 = 4'h7 == io_in[11:8] ? 7'h78 : _GEN_23; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_25 = 4'h8 == io_in[11:8] ? 7'h0 : _GEN_24; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_26 = 4'h9 == io_in[11:8] ? 7'h10 : _GEN_25; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_27 = 4'ha == io_in[11:8] ? 7'h8 : _GEN_26; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_28 = 4'hb == io_in[11:8] ? 7'h3 : _GEN_27; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_29 = 4'hc == io_in[11:8] ? 7'h46 : _GEN_28; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_30 = 4'hd == io_in[11:8] ? 7'h21 : _GEN_29; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_31 = 4'he == io_in[11:8] ? 7'h6 : _GEN_30; // @[SevenSeg.scala 58:20]
  wire [6:0] _GEN_32 = 4'hf == io_in[11:8] ? 7'he : _GEN_31; // @[SevenSeg.scala 58:20]
  wire  _T_12 = 2'h2 == sevAnCounter; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_34 = 4'h1 == io_in[7:4] ? 7'h79 : 7'h40; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_35 = 4'h2 == io_in[7:4] ? 7'h24 : _GEN_34; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_36 = 4'h3 == io_in[7:4] ? 7'h30 : _GEN_35; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_37 = 4'h4 == io_in[7:4] ? 7'h19 : _GEN_36; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_38 = 4'h5 == io_in[7:4] ? 7'h12 : _GEN_37; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_39 = 4'h6 == io_in[7:4] ? 7'h2 : _GEN_38; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_40 = 4'h7 == io_in[7:4] ? 7'h78 : _GEN_39; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_41 = 4'h8 == io_in[7:4] ? 7'h0 : _GEN_40; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_42 = 4'h9 == io_in[7:4] ? 7'h10 : _GEN_41; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_43 = 4'ha == io_in[7:4] ? 7'h8 : _GEN_42; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_44 = 4'hb == io_in[7:4] ? 7'h3 : _GEN_43; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_45 = 4'hc == io_in[7:4] ? 7'h46 : _GEN_44; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_46 = 4'hd == io_in[7:4] ? 7'h21 : _GEN_45; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_47 = 4'he == io_in[7:4] ? 7'h6 : _GEN_46; // @[SevenSeg.scala 62:20]
  wire [6:0] _GEN_48 = 4'hf == io_in[7:4] ? 7'he : _GEN_47; // @[SevenSeg.scala 62:20]
  wire  _T_14 = 2'h3 == sevAnCounter; // @[Conditional.scala 37:30]
  wire [6:0] _GEN_50 = 4'h1 == io_in[3:0] ? 7'h79 : 7'h40; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_51 = 4'h2 == io_in[3:0] ? 7'h24 : _GEN_50; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_52 = 4'h3 == io_in[3:0] ? 7'h30 : _GEN_51; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_53 = 4'h4 == io_in[3:0] ? 7'h19 : _GEN_52; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_54 = 4'h5 == io_in[3:0] ? 7'h12 : _GEN_53; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_55 = 4'h6 == io_in[3:0] ? 7'h2 : _GEN_54; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_56 = 4'h7 == io_in[3:0] ? 7'h78 : _GEN_55; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_57 = 4'h8 == io_in[3:0] ? 7'h0 : _GEN_56; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_58 = 4'h9 == io_in[3:0] ? 7'h10 : _GEN_57; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_59 = 4'ha == io_in[3:0] ? 7'h8 : _GEN_58; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_60 = 4'hb == io_in[3:0] ? 7'h3 : _GEN_59; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_61 = 4'hc == io_in[3:0] ? 7'h46 : _GEN_60; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_62 = 4'hd == io_in[3:0] ? 7'h21 : _GEN_61; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_63 = 4'he == io_in[3:0] ? 7'h6 : _GEN_62; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_64 = 4'hf == io_in[3:0] ? 7'he : _GEN_63; // @[SevenSeg.scala 66:20]
  wire [6:0] _GEN_65 = _T_14 ? _GEN_64 : 7'h0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_66 = _T_14 ? 4'he : 4'h0; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_67 = _T_12 ? _GEN_48 : _GEN_65; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_68 = _T_12 ? 4'hd : _GEN_66; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_69 = _T_10 ? _GEN_32 : _GEN_67; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_70 = _T_10 ? 4'hb : _GEN_68; // @[Conditional.scala 39:67]
  assign io_out_anode = _T_8 ? 4'h7 : _GEN_70; // @[SevenSeg.scala 27:16 SevenSeg.scala 55:20 SevenSeg.scala 59:20 SevenSeg.scala 63:20 SevenSeg.scala 67:20]
  assign io_out_data = _T_8 ? _GEN_16 : _GEN_69; // @[SevenSeg.scala 26:15 SevenSeg.scala 54:20 SevenSeg.scala 58:20 SevenSeg.scala 62:20 SevenSeg.scala 66:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[18:0];
  _RAND_1 = {1{`RANDOM}};
  sevAnCounter = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 19'h0;
    end else if (ticker) begin
      _T <= 19'h0;
    end else begin
      _T <= _T_2;
    end
    if (reset) begin
      sevAnCounter <= 2'h0;
    end else if (ticker) begin
      if (_T_4) begin
        sevAnCounter <= 2'h0;
      end else begin
        sevAnCounter <= _T_6;
      end
    end
  end
endmodule
module Top(
  input         clock,
  input         reset,
  output [15:0] io_blink,
  output [3:0]  io_sev_anode,
  output [6:0]  io_sev_data,
  input         io_ps2_clk,
  input         io_ps2_data,
  input         io_btn
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  mp_clock; // @[Top.scala 18:18]
  wire  mp_reset; // @[Top.scala 18:18]
  wire [31:0] mp_io_dataBus_addr; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_rdData_0; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_rdData_1; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_rdData_2; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_rdData_3; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_wrData_0; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_wrData_1; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_wrData_2; // @[Top.scala 18:18]
  wire [7:0] mp_io_dataBus_wrData_3; // @[Top.scala 18:18]
  wire  mp_io_dataBus_we_0; // @[Top.scala 18:18]
  wire  mp_io_dataBus_we_1; // @[Top.scala 18:18]
  wire  mp_io_dataBus_we_2; // @[Top.scala 18:18]
  wire  mp_io_dataBus_we_3; // @[Top.scala 18:18]
  wire  mp_io_dataBus_w; // @[Top.scala 18:18]
  wire  key_clock; // @[Top.scala 20:19]
  wire  key_reset; // @[Top.scala 20:19]
  wire  key_ps2_clk; // @[Top.scala 20:19]
  wire  key_ps2_data; // @[Top.scala 20:19]
  wire [7:0] key_bus_data; // @[Top.scala 20:19]
  wire [7:0] key_bus_flag; // @[Top.scala 20:19]
  wire  key_bus_clear; // @[Top.scala 20:19]
  wire  ram_clock; // @[Top.scala 24:19]
  wire [31:0] ram_io_addr; // @[Top.scala 24:19]
  wire [7:0] ram_io_rdData_0; // @[Top.scala 24:19]
  wire [7:0] ram_io_rdData_1; // @[Top.scala 24:19]
  wire [7:0] ram_io_rdData_2; // @[Top.scala 24:19]
  wire [7:0] ram_io_rdData_3; // @[Top.scala 24:19]
  wire [7:0] ram_io_wrData_0; // @[Top.scala 24:19]
  wire [7:0] ram_io_wrData_1; // @[Top.scala 24:19]
  wire [7:0] ram_io_wrData_2; // @[Top.scala 24:19]
  wire [7:0] ram_io_wrData_3; // @[Top.scala 24:19]
  wire  ram_io_we_0; // @[Top.scala 24:19]
  wire  ram_io_we_1; // @[Top.scala 24:19]
  wire  ram_io_we_2; // @[Top.scala 24:19]
  wire  ram_io_we_3; // @[Top.scala 24:19]
  wire  ram_io_w; // @[Top.scala 24:19]
  wire  sev_clock; // @[Top.scala 60:19]
  wire  sev_reset; // @[Top.scala 60:19]
  wire [15:0] sev_io_in; // @[Top.scala 60:19]
  wire [3:0] sev_io_out_anode; // @[Top.scala 60:19]
  wire [6:0] sev_io_out_data; // @[Top.scala 60:19]
  reg  _T_2; // @[Top.scala 31:34]
  wire  _T_3 = mp_io_dataBus_w & _T_2; // @[Top.scala 31:24]
  reg  _T_5; // @[Top.scala 35:15]
  wire [7:0] _GEN_4 = _T_5 ? key_bus_flag : ram_io_rdData_0; // @[Top.scala 35:49]
  wire [7:0] _GEN_5 = _T_5 ? 8'h0 : ram_io_rdData_1; // @[Top.scala 35:49]
  wire [7:0] _GEN_6 = _T_5 ? 8'h0 : ram_io_rdData_2; // @[Top.scala 35:49]
  wire [7:0] _GEN_7 = _T_5 ? 8'h0 : ram_io_rdData_3; // @[Top.scala 35:49]
  reg  _T_7; // @[Top.scala 39:15]
  wire [7:0] _GEN_8 = _T_7 ? key_bus_data : _GEN_4; // @[Top.scala 39:49]
  wire [7:0] _GEN_9 = _T_7 ? 8'h0 : _GEN_5; // @[Top.scala 39:49]
  wire [7:0] _GEN_10 = _T_7 ? 8'h0 : _GEN_6; // @[Top.scala 39:49]
  wire [7:0] _GEN_11 = _T_7 ? 8'h0 : _GEN_7; // @[Top.scala 39:49]
  reg  btnReg; // @[Top.scala 45:23]
  wire  _GEN_13 = io_btn | btnReg; // @[Top.scala 46:15]
  reg  _T_9; // @[Top.scala 49:15]
  reg [15:0] blinkReg; // @[Top.scala 55:25]
  reg  _T_11; // @[Top.scala 56:34]
  wire  _T_12 = mp_io_dataBus_w & _T_11; // @[Top.scala 56:24]
  wire [31:0] _T_15 = {mp_io_dataBus_wrData_3,mp_io_dataBus_wrData_2,mp_io_dataBus_wrData_1,mp_io_dataBus_wrData_0}; // @[Cat.scala 29:58]
  RVCore mp ( // @[Top.scala 18:18]
    .clock(mp_clock),
    .reset(mp_reset),
    .io_dataBus_addr(mp_io_dataBus_addr),
    .io_dataBus_rdData_0(mp_io_dataBus_rdData_0),
    .io_dataBus_rdData_1(mp_io_dataBus_rdData_1),
    .io_dataBus_rdData_2(mp_io_dataBus_rdData_2),
    .io_dataBus_rdData_3(mp_io_dataBus_rdData_3),
    .io_dataBus_wrData_0(mp_io_dataBus_wrData_0),
    .io_dataBus_wrData_1(mp_io_dataBus_wrData_1),
    .io_dataBus_wrData_2(mp_io_dataBus_wrData_2),
    .io_dataBus_wrData_3(mp_io_dataBus_wrData_3),
    .io_dataBus_we_0(mp_io_dataBus_we_0),
    .io_dataBus_we_1(mp_io_dataBus_we_1),
    .io_dataBus_we_2(mp_io_dataBus_we_2),
    .io_dataBus_we_3(mp_io_dataBus_we_3),
    .io_dataBus_w(mp_io_dataBus_w)
  );
  PS2 key ( // @[Top.scala 20:19]
    .clock(key_clock),
    .reset(key_reset),
    .ps2_clk(key_ps2_clk),
    .ps2_data(key_ps2_data),
    .bus_data(key_bus_data),
    .bus_flag(key_bus_flag),
    .bus_clear(key_bus_clear)
  );
  RAM ram ( // @[Top.scala 24:19]
    .clock(ram_clock),
    .io_addr(ram_io_addr),
    .io_rdData_0(ram_io_rdData_0),
    .io_rdData_1(ram_io_rdData_1),
    .io_rdData_2(ram_io_rdData_2),
    .io_rdData_3(ram_io_rdData_3),
    .io_wrData_0(ram_io_wrData_0),
    .io_wrData_1(ram_io_wrData_1),
    .io_wrData_2(ram_io_wrData_2),
    .io_wrData_3(ram_io_wrData_3),
    .io_we_0(ram_io_we_0),
    .io_we_1(ram_io_we_1),
    .io_we_2(ram_io_we_2),
    .io_we_3(ram_io_we_3),
    .io_w(ram_io_w)
  );
  SevenSeg sev ( // @[Top.scala 60:19]
    .clock(sev_clock),
    .reset(sev_reset),
    .io_in(sev_io_in),
    .io_out_anode(sev_io_out_anode),
    .io_out_data(sev_io_out_data)
  );
  assign io_blink = blinkReg; // @[Top.scala 59:12]
  assign io_sev_anode = sev_io_out_anode; // @[Top.scala 61:14]
  assign io_sev_data = sev_io_out_data; // @[Top.scala 61:14]
  assign mp_clock = clock;
  assign mp_reset = reset;
  assign mp_io_dataBus_rdData_0 = _T_9 ? {{7'd0}, btnReg} : _GEN_8; // @[Top.scala 25:24 Top.scala 36:26 Top.scala 37:29 Top.scala 40:26 Top.scala 41:29 Top.scala 50:26 Top.scala 51:29]
  assign mp_io_dataBus_rdData_1 = _T_9 ? 8'h0 : _GEN_9; // @[Top.scala 25:24 Top.scala 36:26 Top.scala 40:26 Top.scala 50:26]
  assign mp_io_dataBus_rdData_2 = _T_9 ? 8'h0 : _GEN_10; // @[Top.scala 25:24 Top.scala 36:26 Top.scala 40:26 Top.scala 50:26]
  assign mp_io_dataBus_rdData_3 = _T_9 ? 8'h0 : _GEN_11; // @[Top.scala 25:24 Top.scala 36:26 Top.scala 40:26 Top.scala 50:26]
  assign key_clock = clock;
  assign key_reset = reset;
  assign key_ps2_clk = io_ps2_clk; // @[Top.scala 21:11]
  assign key_ps2_data = io_ps2_data; // @[Top.scala 21:11]
  assign key_bus_clear = _T_7; // @[Top.scala 22:17 Top.scala 42:19]
  assign ram_clock = clock;
  assign ram_io_addr = mp_io_dataBus_addr; // @[Top.scala 27:15]
  assign ram_io_wrData_0 = mp_io_dataBus_wrData_0; // @[Top.scala 28:17]
  assign ram_io_wrData_1 = mp_io_dataBus_wrData_1; // @[Top.scala 28:17]
  assign ram_io_wrData_2 = mp_io_dataBus_wrData_2; // @[Top.scala 28:17]
  assign ram_io_wrData_3 = mp_io_dataBus_wrData_3; // @[Top.scala 28:17]
  assign ram_io_we_0 = _T_3 & mp_io_dataBus_we_0; // @[Top.scala 29:13 Top.scala 32:15]
  assign ram_io_we_1 = _T_3 & mp_io_dataBus_we_1; // @[Top.scala 29:13 Top.scala 32:15]
  assign ram_io_we_2 = _T_3 & mp_io_dataBus_we_2; // @[Top.scala 29:13 Top.scala 32:15]
  assign ram_io_we_3 = _T_3 & mp_io_dataBus_we_3; // @[Top.scala 29:13 Top.scala 32:15]
  assign ram_io_w = mp_io_dataBus_w; // @[Top.scala 30:12]
  assign sev_clock = clock;
  assign sev_reset = reset;
  assign sev_io_in = blinkReg; // @[Top.scala 62:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_7 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  btnReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_9 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  blinkReg = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  _T_11 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_2 <= mp_io_dataBus_addr <= 32'h1000;
    _T_5 <= mp_io_dataBus_addr == 32'h2100;
    _T_7 <= mp_io_dataBus_addr == 32'h2200;
    if (reset) begin
      btnReg <= 1'h0;
    end else if (_T_9) begin
      btnReg <= 1'h0;
    end else begin
      btnReg <= _GEN_13;
    end
    _T_9 <= mp_io_dataBus_addr == 32'h2300;
    if (reset) begin
      blinkReg <= 16'h0;
    end else if (_T_12) begin
      blinkReg <= _T_15[15:0];
    end
    _T_11 <= mp_io_dataBus_addr == 32'h2000;
  end
endmodule
