module IF(
  input         clock,
  input         reset,
  input  [31:0] in_pcNext,
  input         in_branch,
  output [31:0] out_pc,
  output [31:0] out_instr,
  output [31:0] instrBus_pc,
  input  [31:0] instrBus_instr,
  input         ctrl_pcEn
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[IF.scala 19:19]
  wire [31:0] _T_3 = pc + 32'h4; // @[IF.scala 52:14]
  assign out_pc = pc; // @[IF.scala 47:10]
  assign out_instr = instrBus_instr; // @[IF.scala 45:13]
  assign instrBus_pc = pc; // @[IF.scala 24:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h0;
    end else if (ctrl_pcEn) begin
      if (in_branch) begin
        pc <= in_pcNext;
      end else begin
        pc <= _T_3;
      end
    end
  end
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_registerS1Index,
  input  [4:0]  io_registerS2Index,
  input  [4:0]  io_registerWIndex,
  input  [31:0] io_registerWData,
  input         io_writeEn,
  output [31:0] io_registerS1Data,
  output [31:0] io_registerS2Data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regFile_1; // @[RegFile.scala 17:24]
  reg [31:0] regFile_2; // @[RegFile.scala 17:24]
  reg [31:0] regFile_3; // @[RegFile.scala 17:24]
  reg [31:0] regFile_4; // @[RegFile.scala 17:24]
  reg [31:0] regFile_5; // @[RegFile.scala 17:24]
  reg [31:0] regFile_6; // @[RegFile.scala 17:24]
  reg [31:0] regFile_7; // @[RegFile.scala 17:24]
  reg [31:0] regFile_8; // @[RegFile.scala 17:24]
  reg [31:0] regFile_9; // @[RegFile.scala 17:24]
  reg [31:0] regFile_10; // @[RegFile.scala 17:24]
  reg [31:0] regFile_11; // @[RegFile.scala 17:24]
  reg [31:0] regFile_12; // @[RegFile.scala 17:24]
  reg [31:0] regFile_13; // @[RegFile.scala 17:24]
  reg [31:0] regFile_14; // @[RegFile.scala 17:24]
  reg [31:0] regFile_15; // @[RegFile.scala 17:24]
  reg [31:0] regFile_16; // @[RegFile.scala 17:24]
  reg [31:0] regFile_17; // @[RegFile.scala 17:24]
  reg [31:0] regFile_18; // @[RegFile.scala 17:24]
  reg [31:0] regFile_19; // @[RegFile.scala 17:24]
  reg [31:0] regFile_20; // @[RegFile.scala 17:24]
  reg [31:0] regFile_21; // @[RegFile.scala 17:24]
  reg [31:0] regFile_22; // @[RegFile.scala 17:24]
  reg [31:0] regFile_23; // @[RegFile.scala 17:24]
  reg [31:0] regFile_24; // @[RegFile.scala 17:24]
  reg [31:0] regFile_25; // @[RegFile.scala 17:24]
  reg [31:0] regFile_26; // @[RegFile.scala 17:24]
  reg [31:0] regFile_27; // @[RegFile.scala 17:24]
  reg [31:0] regFile_28; // @[RegFile.scala 17:24]
  reg [31:0] regFile_29; // @[RegFile.scala 17:24]
  reg [31:0] regFile_30; // @[RegFile.scala 17:24]
  reg [31:0] regFile_31; // @[RegFile.scala 17:24]
  wire [31:0] _GEN_65 = 5'h1 == io_registerS1Index ? $signed(regFile_1) : $signed(32'sh0); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_66 = 5'h2 == io_registerS1Index ? $signed(regFile_2) : $signed(_GEN_65); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_67 = 5'h3 == io_registerS1Index ? $signed(regFile_3) : $signed(_GEN_66); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_68 = 5'h4 == io_registerS1Index ? $signed(regFile_4) : $signed(_GEN_67); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_69 = 5'h5 == io_registerS1Index ? $signed(regFile_5) : $signed(_GEN_68); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_70 = 5'h6 == io_registerS1Index ? $signed(regFile_6) : $signed(_GEN_69); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_71 = 5'h7 == io_registerS1Index ? $signed(regFile_7) : $signed(_GEN_70); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_72 = 5'h8 == io_registerS1Index ? $signed(regFile_8) : $signed(_GEN_71); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_73 = 5'h9 == io_registerS1Index ? $signed(regFile_9) : $signed(_GEN_72); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_74 = 5'ha == io_registerS1Index ? $signed(regFile_10) : $signed(_GEN_73); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_75 = 5'hb == io_registerS1Index ? $signed(regFile_11) : $signed(_GEN_74); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_76 = 5'hc == io_registerS1Index ? $signed(regFile_12) : $signed(_GEN_75); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_77 = 5'hd == io_registerS1Index ? $signed(regFile_13) : $signed(_GEN_76); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_78 = 5'he == io_registerS1Index ? $signed(regFile_14) : $signed(_GEN_77); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_79 = 5'hf == io_registerS1Index ? $signed(regFile_15) : $signed(_GEN_78); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_80 = 5'h10 == io_registerS1Index ? $signed(regFile_16) : $signed(_GEN_79); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_81 = 5'h11 == io_registerS1Index ? $signed(regFile_17) : $signed(_GEN_80); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_82 = 5'h12 == io_registerS1Index ? $signed(regFile_18) : $signed(_GEN_81); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_83 = 5'h13 == io_registerS1Index ? $signed(regFile_19) : $signed(_GEN_82); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_84 = 5'h14 == io_registerS1Index ? $signed(regFile_20) : $signed(_GEN_83); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_85 = 5'h15 == io_registerS1Index ? $signed(regFile_21) : $signed(_GEN_84); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_86 = 5'h16 == io_registerS1Index ? $signed(regFile_22) : $signed(_GEN_85); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_87 = 5'h17 == io_registerS1Index ? $signed(regFile_23) : $signed(_GEN_86); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_88 = 5'h18 == io_registerS1Index ? $signed(regFile_24) : $signed(_GEN_87); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_89 = 5'h19 == io_registerS1Index ? $signed(regFile_25) : $signed(_GEN_88); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_90 = 5'h1a == io_registerS1Index ? $signed(regFile_26) : $signed(_GEN_89); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_91 = 5'h1b == io_registerS1Index ? $signed(regFile_27) : $signed(_GEN_90); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_92 = 5'h1c == io_registerS1Index ? $signed(regFile_28) : $signed(_GEN_91); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_93 = 5'h1d == io_registerS1Index ? $signed(regFile_29) : $signed(_GEN_92); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_94 = 5'h1e == io_registerS1Index ? $signed(regFile_30) : $signed(_GEN_93); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_95 = 5'h1f == io_registerS1Index ? $signed(regFile_31) : $signed(_GEN_94); // @[RegFile.scala 24:21]
  wire [31:0] _GEN_97 = 5'h1 == io_registerS2Index ? $signed(regFile_1) : $signed(32'sh0); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_98 = 5'h2 == io_registerS2Index ? $signed(regFile_2) : $signed(_GEN_97); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_99 = 5'h3 == io_registerS2Index ? $signed(regFile_3) : $signed(_GEN_98); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_100 = 5'h4 == io_registerS2Index ? $signed(regFile_4) : $signed(_GEN_99); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_101 = 5'h5 == io_registerS2Index ? $signed(regFile_5) : $signed(_GEN_100); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_102 = 5'h6 == io_registerS2Index ? $signed(regFile_6) : $signed(_GEN_101); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_103 = 5'h7 == io_registerS2Index ? $signed(regFile_7) : $signed(_GEN_102); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_104 = 5'h8 == io_registerS2Index ? $signed(regFile_8) : $signed(_GEN_103); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_105 = 5'h9 == io_registerS2Index ? $signed(regFile_9) : $signed(_GEN_104); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_106 = 5'ha == io_registerS2Index ? $signed(regFile_10) : $signed(_GEN_105); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_107 = 5'hb == io_registerS2Index ? $signed(regFile_11) : $signed(_GEN_106); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_108 = 5'hc == io_registerS2Index ? $signed(regFile_12) : $signed(_GEN_107); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_109 = 5'hd == io_registerS2Index ? $signed(regFile_13) : $signed(_GEN_108); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_110 = 5'he == io_registerS2Index ? $signed(regFile_14) : $signed(_GEN_109); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_111 = 5'hf == io_registerS2Index ? $signed(regFile_15) : $signed(_GEN_110); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_112 = 5'h10 == io_registerS2Index ? $signed(regFile_16) : $signed(_GEN_111); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_113 = 5'h11 == io_registerS2Index ? $signed(regFile_17) : $signed(_GEN_112); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_114 = 5'h12 == io_registerS2Index ? $signed(regFile_18) : $signed(_GEN_113); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_115 = 5'h13 == io_registerS2Index ? $signed(regFile_19) : $signed(_GEN_114); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_116 = 5'h14 == io_registerS2Index ? $signed(regFile_20) : $signed(_GEN_115); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_117 = 5'h15 == io_registerS2Index ? $signed(regFile_21) : $signed(_GEN_116); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_118 = 5'h16 == io_registerS2Index ? $signed(regFile_22) : $signed(_GEN_117); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_119 = 5'h17 == io_registerS2Index ? $signed(regFile_23) : $signed(_GEN_118); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_120 = 5'h18 == io_registerS2Index ? $signed(regFile_24) : $signed(_GEN_119); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_121 = 5'h19 == io_registerS2Index ? $signed(regFile_25) : $signed(_GEN_120); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_122 = 5'h1a == io_registerS2Index ? $signed(regFile_26) : $signed(_GEN_121); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_123 = 5'h1b == io_registerS2Index ? $signed(regFile_27) : $signed(_GEN_122); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_124 = 5'h1c == io_registerS2Index ? $signed(regFile_28) : $signed(_GEN_123); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_125 = 5'h1d == io_registerS2Index ? $signed(regFile_29) : $signed(_GEN_124); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_126 = 5'h1e == io_registerS2Index ? $signed(regFile_30) : $signed(_GEN_125); // @[RegFile.scala 25:21]
  wire [31:0] _GEN_127 = 5'h1f == io_registerS2Index ? $signed(regFile_31) : $signed(_GEN_126); // @[RegFile.scala 25:21]
  wire  _T_1 = io_registerS1Index == io_registerWIndex; // @[RegFile.scala 27:27]
  wire  _T_2 = io_registerS1Index != 5'h0; // @[RegFile.scala 27:71]
  wire  _T_3 = _T_1 & _T_2; // @[RegFile.scala 27:49]
  wire  _T_4 = _T_3 & io_writeEn; // @[RegFile.scala 27:79]
  wire  _T_5 = io_registerS2Index == io_registerWIndex; // @[RegFile.scala 30:27]
  wire  _T_6 = io_registerS2Index != 5'h0; // @[RegFile.scala 30:71]
  wire  _T_7 = _T_5 & _T_6; // @[RegFile.scala 30:49]
  wire  _T_8 = _T_7 & io_writeEn; // @[RegFile.scala 30:79]
  assign io_registerS1Data = _T_4 ? $signed(io_registerWData) : $signed(_GEN_95); // @[RegFile.scala 24:21 RegFile.scala 28:23]
  assign io_registerS2Data = _T_8 ? $signed(io_registerWData) : $signed(_GEN_127); // @[RegFile.scala 25:21 RegFile.scala 31:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regFile_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regFile_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regFile_3 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regFile_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regFile_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regFile_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regFile_7 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regFile_8 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regFile_9 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regFile_10 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regFile_11 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regFile_12 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regFile_13 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regFile_14 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regFile_15 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regFile_16 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regFile_17 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regFile_18 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regFile_19 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regFile_20 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regFile_21 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regFile_22 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regFile_23 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regFile_24 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regFile_25 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regFile_26 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regFile_27 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regFile_28 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regFile_29 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regFile_30 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regFile_31 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regFile_1 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1 == io_registerWIndex) begin
        regFile_1 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_2 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h2 == io_registerWIndex) begin
        regFile_2 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_3 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h3 == io_registerWIndex) begin
        regFile_3 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_4 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h4 == io_registerWIndex) begin
        regFile_4 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_5 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h5 == io_registerWIndex) begin
        regFile_5 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_6 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h6 == io_registerWIndex) begin
        regFile_6 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_7 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h7 == io_registerWIndex) begin
        regFile_7 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_8 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h8 == io_registerWIndex) begin
        regFile_8 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_9 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h9 == io_registerWIndex) begin
        regFile_9 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_10 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'ha == io_registerWIndex) begin
        regFile_10 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_11 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hb == io_registerWIndex) begin
        regFile_11 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_12 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hc == io_registerWIndex) begin
        regFile_12 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_13 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hd == io_registerWIndex) begin
        regFile_13 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_14 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'he == io_registerWIndex) begin
        regFile_14 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_15 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'hf == io_registerWIndex) begin
        regFile_15 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_16 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h10 == io_registerWIndex) begin
        regFile_16 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_17 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h11 == io_registerWIndex) begin
        regFile_17 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_18 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h12 == io_registerWIndex) begin
        regFile_18 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_19 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h13 == io_registerWIndex) begin
        regFile_19 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_20 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h14 == io_registerWIndex) begin
        regFile_20 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_21 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h15 == io_registerWIndex) begin
        regFile_21 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_22 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h16 == io_registerWIndex) begin
        regFile_22 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_23 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h17 == io_registerWIndex) begin
        regFile_23 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_24 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h18 == io_registerWIndex) begin
        regFile_24 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_25 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h19 == io_registerWIndex) begin
        regFile_25 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_26 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1a == io_registerWIndex) begin
        regFile_26 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_27 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1b == io_registerWIndex) begin
        regFile_27 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_28 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1c == io_registerWIndex) begin
        regFile_28 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_29 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1d == io_registerWIndex) begin
        regFile_29 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_30 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1e == io_registerWIndex) begin
        regFile_30 <= io_registerWData;
      end
    end
    if (reset) begin
      regFile_31 <= 32'sh0;
    end else if (io_writeEn) begin
      if (5'h1f == io_registerWIndex) begin
        regFile_31 <= io_registerWData;
      end
    end
  end
endmodule
module ImmGen(
  input  [31:0] io_instruction,
  output [31:0] io_immediate
);
  wire [2:0] funct3 = io_instruction[14:12]; // @[ImmGen.scala 13:30]
  wire [11:0] Itype = io_instruction[31:20]; // @[ImmGen.scala 19:29]
  wire [9:0] _T_45 = {io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31]}; // @[ImmGen.scala 21:71]
  wire [31:0] _T_57 = {_T_45,_T_45,Itype}; // @[ImmGen.scala 21:88]
  wire  _T_58 = funct3 == 3'h2; // @[ImmGen.scala 22:15]
  wire  _T_59 = funct3 == 3'h3; // @[ImmGen.scala 22:33]
  wire  _T_60 = _T_58 | _T_59; // @[ImmGen.scala 22:23]
  wire [11:0] _T_61 = io_instruction[31:20]; // @[ImmGen.scala 23:33]
  wire [31:0] _GEN_0 = _T_60 ? $signed({{20{_T_61[11]}},_T_61}) : $signed(_T_57); // @[ImmGen.scala 22:42]
  wire  _T_63 = 7'h37 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [31:0] _T_64 = {io_instruction[31:12],12'h0}; // @[ImmGen.scala 29:35]
  wire  _T_65 = 7'h17 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire  _T_67 = 7'h6f == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [30:0] _T_90 = {_T_45,io_instruction[31],io_instruction[19:12],io_instruction[20],io_instruction[30:22],2'h0}; // @[ImmGen.scala 35:103]
  wire  _T_91 = 7'h23 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [31:0] _T_133 = {_T_45,_T_45,io_instruction[31:25],io_instruction[11:7]}; // @[ImmGen.scala 38:92]
  wire  _T_134 = 7'h63 == io_instruction[6:0]; // @[Conditional.scala 37:30]
  wire [8:0] _T_161 = {io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31]}; // @[ImmGen.scala 41:75]
  wire [17:0] _T_170 = {io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],io_instruction[31],_T_161}; // @[ImmGen.scala 41:75]
  wire [30:0] _T_173 = {_T_170,io_instruction[31],io_instruction[7],io_instruction[30:25],io_instruction[11:8],1'h0}; // @[ImmGen.scala 41:103]
  wire [31:0] _GEN_1 = _T_134 ? $signed({{1{_T_173[30]}},_T_173}) : $signed(_GEN_0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_91 ? $signed(_T_133) : $signed(_GEN_1); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_3 = _T_67 ? $signed({{1{_T_90[30]}},_T_90}) : $signed(_GEN_2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_4 = _T_65 ? $signed(_T_64) : $signed(_GEN_3); // @[Conditional.scala 39:67]
  assign io_immediate = _T_63 ? $signed(_T_64) : $signed(_GEN_4); // @[ImmGen.scala 21:16 ImmGen.scala 23:18 ImmGen.scala 29:20 ImmGen.scala 32:20 ImmGen.scala 35:20 ImmGen.scala 38:20 ImmGen.scala 41:20]
endmodule
module ID(
  input         clock,
  input         reset,
  input  [31:0] in_pc,
  input  [31:0] in_instr,
  output [31:0] out_pc,
  output [31:0] out_imm,
  output [31:0] out_regOp1,
  output [31:0] out_regOp2,
  output [4:0]  out_rs1,
  output [4:0]  out_rs2,
  output [4:0]  out_rd,
  output [3:0]  out_aluOp,
  output [1:0]  out_aluSrc1,
  output [1:0]  out_aluSrc2,
  output        out_brSrc,
  output        out_pcSrc,
  output        out_wb,
  output        out_wbSrc,
  output [3:0]  out_mem,
  output        out_jump,
  output [2:0]  out_funct3,
  input  [4:0]  wb_rd,
  input  [31:0] wb_res,
  input         wb_wb,
  input         ctrl_flushID,
  output [31:0] ctrl_instr
);
  wire  regFile_clock; // @[ID.scala 22:23]
  wire  regFile_reset; // @[ID.scala 22:23]
  wire [4:0] regFile_io_registerS1Index; // @[ID.scala 22:23]
  wire [4:0] regFile_io_registerS2Index; // @[ID.scala 22:23]
  wire [4:0] regFile_io_registerWIndex; // @[ID.scala 22:23]
  wire [31:0] regFile_io_registerWData; // @[ID.scala 22:23]
  wire  regFile_io_writeEn; // @[ID.scala 22:23]
  wire [31:0] regFile_io_registerS1Data; // @[ID.scala 22:23]
  wire [31:0] regFile_io_registerS2Data; // @[ID.scala 22:23]
  wire [31:0] immGen_io_instruction; // @[ID.scala 24:22]
  wire [31:0] immGen_io_immediate; // @[ID.scala 24:22]
  wire [6:0] opcode = in_instr[6:0]; // @[ID.scala 26:24]
  wire [2:0] funct3 = in_instr[14:12]; // @[ID.scala 27:24]
  wire  _T_1 = 7'h3 == opcode; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h0 == funct3; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h4 == funct3; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h1 == funct3; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h5 == funct3; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h2 == funct3; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_0 = _T_6 ? 3'h7 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1 = _T_5 ? 3'h2 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_4 ? 3'h6 : _GEN_1; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_3 = _T_3 ? 3'h1 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_2 ? 3'h5 : _GEN_3; // @[Conditional.scala 40:58]
  wire  _T_7 = 7'h23 == opcode; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_5 = _T_6 ? 4'hb : 4'h0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_6 = _T_4 ? 4'ha : _GEN_5; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_7 = _T_2 ? 4'h9 : _GEN_6; // @[Conditional.scala 40:58]
  wire  _T_11 = 7'h13 == opcode; // @[Conditional.scala 37:30]
  wire  _T_15 = 3'h3 == funct3; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_8 = in_instr[30] ? 4'h4 : 4'h3; // @[ID.scala 119:30]
  wire  _T_19 = 3'h6 == funct3; // @[Conditional.scala 37:30]
  wire  _T_20 = 3'h7 == funct3; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_9 = _T_20 ? 4'h5 : 4'h0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_10 = _T_19 ? 4'h6 : _GEN_9; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_11 = _T_5 ? _GEN_8 : _GEN_10; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_12 = _T_3 ? 4'h7 : _GEN_11; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_13 = _T_15 ? 4'h8 : _GEN_12; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_14 = _T_6 ? 4'h8 : _GEN_13; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_15 = _T_4 ? 4'h2 : _GEN_14; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_16 = _T_2 ? 4'h0 : _GEN_15; // @[Conditional.scala 40:58]
  wire  _T_21 = 7'h33 == opcode; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_17 = in_instr[30] ? 4'h1 : 4'h0; // @[ID.scala 136:30]
  wire [3:0] _GEN_26 = _T_2 ? _GEN_17 : _GEN_15; // @[Conditional.scala 40:58]
  wire  _T_32 = 7'h17 == opcode; // @[Conditional.scala 37:30]
  wire  _T_33 = 7'h37 == opcode; // @[Conditional.scala 37:30]
  wire  _T_34 = 7'h63 == opcode; // @[Conditional.scala 37:30]
  wire  _T_35 = 7'h6f == opcode; // @[Conditional.scala 37:30]
  wire  _T_36 = 7'h67 == opcode; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_28 = _T_36 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_35 | _T_36; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_30 = _T_35 ? 2'h1 : _GEN_28; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_31 = _T_35 ? 2'h2 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_32 = _T_35 ? 1'h0 : _T_36; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_34 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_34 | _GEN_29; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_35 = _T_34 ? 2'h0 : _GEN_30; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_36 = _T_34 ? 2'h0 : _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_34 ? 1'h0 : _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_33 | _GEN_33; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_39 = _T_33 ? 2'h2 : _GEN_35; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_40 = _T_33 ? 2'h1 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_33 ? 1'h0 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_33 ? 1'h0 : _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_32 | _GEN_38; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_44 = _T_32 ? 2'h1 : _GEN_39; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_45 = _T_32 ? 2'h1 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_46 = _T_32 ? 1'h0 : _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_32 ? 1'h0 : _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_21 | _GEN_43; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_49 = _T_21 ? _GEN_26 : 4'h0; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_50 = _T_21 ? 2'h0 : _GEN_44; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_51 = _T_21 ? 2'h0 : _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_21 ? 1'h0 : _GEN_46; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_21 ? 1'h0 : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_11 | _GEN_48; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_55 = _T_11 ? 2'h1 : _GEN_51; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_56 = _T_11 ? _GEN_16 : _GEN_49; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_57 = _T_11 ? 2'h0 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_11 ? 1'h0 : _GEN_52; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_11 ? 1'h0 : _GEN_53; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_60 = _T_7 ? 2'h1 : _GEN_55; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_61 = _T_7 ? _GEN_7 : 4'h0; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_7 ? 1'h0 : _GEN_54; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_63 = _T_7 ? 4'h0 : _GEN_56; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_64 = _T_7 ? 2'h0 : _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_7 ? 1'h0 : _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_7 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_1 | _GEN_62; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_70 = _T_1 ? {{1'd0}, _GEN_4} : _GEN_61; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_71 = _T_1 ? 4'h0 : _GEN_63; // @[Conditional.scala 40:58]
  wire  _GEN_73 = _T_1 ? 1'h0 : _GEN_65; // @[Conditional.scala 40:58]
  RegFile regFile ( // @[ID.scala 22:23]
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_registerS1Index(regFile_io_registerS1Index),
    .io_registerS2Index(regFile_io_registerS2Index),
    .io_registerWIndex(regFile_io_registerWIndex),
    .io_registerWData(regFile_io_registerWData),
    .io_writeEn(regFile_io_writeEn),
    .io_registerS1Data(regFile_io_registerS1Data),
    .io_registerS2Data(regFile_io_registerS2Data)
  );
  ImmGen immGen ( // @[ID.scala 24:22]
    .io_instruction(immGen_io_instruction),
    .io_immediate(immGen_io_immediate)
  );
  assign out_pc = in_pc; // @[ID.scala 51:10]
  assign out_imm = immGen_io_immediate; // @[ID.scala 46:11]
  assign out_regOp1 = regFile_io_registerS1Data; // @[ID.scala 38:14]
  assign out_regOp2 = regFile_io_registerS2Data; // @[ID.scala 39:14]
  assign out_rs1 = in_instr[19:15]; // @[ID.scala 48:11]
  assign out_rs2 = in_instr[24:20]; // @[ID.scala 49:11]
  assign out_rd = in_instr[11:7]; // @[ID.scala 50:10]
  assign out_aluOp = ctrl_flushID ? 4'h0 : _GEN_71; // @[ID.scala 55:13 ID.scala 103:21 ID.scala 106:21 ID.scala 109:21 ID.scala 112:21 ID.scala 115:21 ID.scala 118:21 ID.scala 120:23 ID.scala 124:21 ID.scala 127:21 ID.scala 135:21 ID.scala 137:23 ID.scala 141:21 ID.scala 144:21 ID.scala 147:21 ID.scala 150:21 ID.scala 153:21 ID.scala 155:23 ID.scala 159:21 ID.scala 162:21 ID.scala 198:15]
  assign out_aluSrc1 = _T_1 ? 2'h0 : _GEN_64; // @[ID.scala 53:15 ID.scala 168:19 ID.scala 173:19 ID.scala 182:19 ID.scala 189:19]
  assign out_aluSrc2 = _T_1 ? 2'h1 : _GEN_60; // @[ID.scala 54:15 ID.scala 64:19 ID.scala 85:19 ID.scala 100:19 ID.scala 169:19 ID.scala 174:19 ID.scala 183:19 ID.scala 190:19]
  assign out_brSrc = _T_1 ? 1'h0 : _GEN_66; // @[ID.scala 59:13 ID.scala 188:17]
  assign out_pcSrc = ctrl_flushID ? 1'h0 : _GEN_73; // @[ID.scala 57:13 ID.scala 178:17 ID.scala 184:17 ID.scala 191:17 ID.scala 201:15]
  assign out_wb = ctrl_flushID ? 1'h0 : _GEN_67; // @[ID.scala 52:10 ID.scala 63:14 ID.scala 99:14 ID.scala 132:14 ID.scala 167:14 ID.scala 172:14 ID.scala 177:14 ID.scala 181:14 ID.scala 187:14 ID.scala 197:12]
  assign out_wbSrc = ctrl_flushID ? 1'h0 : _T_1; // @[ID.scala 58:13 ID.scala 65:17 ID.scala 200:15]
  assign out_mem = ctrl_flushID ? 4'h0 : _GEN_70; // @[ID.scala 56:11 ID.scala 68:19 ID.scala 71:19 ID.scala 74:19 ID.scala 77:19 ID.scala 80:19 ID.scala 88:19 ID.scala 91:19 ID.scala 94:19 ID.scala 199:13]
  assign out_jump = opcode[2]; // @[ID.scala 32:12]
  assign out_funct3 = in_instr[14:12]; // @[ID.scala 33:14]
  assign ctrl_instr = in_instr; // @[ID.scala 195:14]
  assign regFile_clock = clock;
  assign regFile_reset = reset;
  assign regFile_io_registerS1Index = in_instr[19:15]; // @[ID.scala 36:30]
  assign regFile_io_registerS2Index = in_instr[24:20]; // @[ID.scala 37:30]
  assign regFile_io_registerWIndex = wb_rd; // @[ID.scala 41:29]
  assign regFile_io_registerWData = wb_res; // @[ID.scala 42:28]
  assign regFile_io_writeEn = wb_wb; // @[ID.scala 43:22]
  assign immGen_io_instruction = in_instr; // @[ID.scala 45:25]
endmodule
module ALU(
  input  [31:0] io_source1,
  input  [31:0] io_source2,
  input  [3:0]  io_operation,
  output [31:0] io_output
);
  wire [31:0] _T_2 = $signed(io_source1) + $signed(io_source2); // @[ALU.scala 19:27]
  wire  _T_3 = 4'h1 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_6 = $signed(io_source1) - $signed(io_source2); // @[ALU.scala 23:31]
  wire  _T_7 = 4'h2 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_8 = io_source1; // @[ALU.scala 26:32]
  wire [62:0] _GEN_8 = {{31'd0}, _T_8}; // @[ALU.scala 26:39]
  wire [62:0] _T_11 = _GEN_8 << io_source2[4:0]; // @[ALU.scala 26:67]
  wire  _T_12 = 4'h3 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_16 = io_source1 >> io_source2[4:0]; // @[ALU.scala 29:67]
  wire  _T_17 = 4'h4 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_19 = $signed(io_source1) >>> io_source2[4:0]; // @[ALU.scala 32:32]
  wire  _T_20 = 4'h6 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_22 = $signed(io_source1) | $signed(io_source2); // @[ALU.scala 35:31]
  wire  _T_23 = 4'h5 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_25 = $signed(io_source1) & $signed(io_source2); // @[ALU.scala 38:31]
  wire  _T_26 = 4'h7 == io_operation; // @[Conditional.scala 37:30]
  wire [31:0] _T_28 = $signed(io_source1) ^ $signed(io_source2); // @[ALU.scala 41:31]
  wire  _T_29 = 4'h8 == io_operation; // @[Conditional.scala 37:30]
  wire  _T_31 = $signed(io_source1) < $signed(io_source2); // @[ALU.scala 44:52]
  wire [31:0] _GEN_0 = _T_29 ? $signed({32{_T_31}}) : $signed(_T_2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1 = _T_26 ? $signed(_T_28) : $signed(_GEN_0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_23 ? $signed(_T_25) : $signed(_GEN_1); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_3 = _T_20 ? $signed(_T_22) : $signed(_GEN_2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_4 = _T_17 ? $signed(_T_19) : $signed(_GEN_3); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5 = _T_12 ? $signed(_T_16) : $signed(_GEN_4); // @[Conditional.scala 39:67]
  wire [62:0] _GEN_6 = _T_7 ? $signed(_T_11) : $signed({{31{_GEN_5[31]}},_GEN_5}); // @[Conditional.scala 39:67]
  wire [62:0] _GEN_7 = _T_3 ? $signed({{31{_T_6[31]}},_T_6}) : $signed(_GEN_6); // @[Conditional.scala 40:58]
  assign io_output = _GEN_7[31:0]; // @[ALU.scala 19:13 ALU.scala 23:17 ALU.scala 26:17 ALU.scala 29:17 ALU.scala 32:17 ALU.scala 35:17 ALU.scala 38:17 ALU.scala 41:17 ALU.scala 44:17]
endmodule
module BranchControl(
  input  [2:0]  io_funct3,
  input  [31:0] io_registerS1,
  input  [31:0] io_registerS2,
  input         io_jump,
  output        io_takeBranch
);
  wire  equal = $signed(io_registerS1) == $signed(io_registerS2); // @[BranchControl.scala 15:29]
  wire  lessThan = $signed(io_registerS1) < $signed(io_registerS2); // @[BranchControl.scala 16:32]
  wire  lessThanU = io_registerS1 < io_registerS2; // @[BranchControl.scala 17:42]
  wire  _T_2 = 3'h0 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h1 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_4 = ~equal; // @[BranchControl.scala 26:24]
  wire  _T_5 = 3'h4 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h5 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_7 = ~lessThan; // @[BranchControl.scala 32:24]
  wire  _T_8 = 3'h6 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h7 == io_funct3; // @[Conditional.scala 37:30]
  wire  _T_10 = ~lessThanU; // @[BranchControl.scala 38:24]
  wire  _GEN_0 = _T_9 & _T_10; // @[Conditional.scala 39:67]
  wire  _GEN_1 = _T_8 ? lessThanU : _GEN_0; // @[Conditional.scala 39:67]
  wire  _GEN_2 = _T_6 ? _T_7 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_5 ? lessThan : _GEN_2; // @[Conditional.scala 39:67]
  wire  _GEN_4 = _T_3 ? _T_4 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_2 ? equal : _GEN_4; // @[Conditional.scala 40:58]
  assign io_takeBranch = io_jump | _GEN_5; // @[BranchControl.scala 19:17 BranchControl.scala 23:21 BranchControl.scala 26:21 BranchControl.scala 29:21 BranchControl.scala 32:21 BranchControl.scala 35:21 BranchControl.scala 38:21 BranchControl.scala 42:19]
endmodule
module EX(
  input  [31:0] in_pc,
  input  [31:0] in_imm,
  input  [31:0] in_regOp1,
  input  [31:0] in_regOp2,
  input  [4:0]  in_rs1,
  input  [4:0]  in_rs2,
  input  [4:0]  in_rd,
  input  [3:0]  in_aluOp,
  input  [1:0]  in_aluSrc1,
  input  [1:0]  in_aluSrc2,
  input         in_brSrc,
  input         in_pcSrc,
  input         in_wb,
  input         in_wbSrc,
  input  [3:0]  in_mem,
  input         in_jump,
  input  [2:0]  in_funct3,
  output [31:0] out_aluRes,
  output [4:0]  out_rd,
  output        out_wb,
  output        out_wbSrc,
  output [3:0]  out_mem,
  output [4:0]  ctrl_rs1,
  output [4:0]  ctrl_rs2,
  output [4:0]  ctrl_rd,
  input  [31:0] ctrl_fwdA,
  input  [31:0] ctrl_fwdB,
  input         ctrl_fwdA_en,
  input         ctrl_fwdB_en,
  output [31:0] ctrl_branchOut_pcNext,
  output        ctrl_branchOut_branch,
  output [1:0]  sysBusMaster_cmd,
  output [31:0] sysBusMaster_addr,
  output [31:0] sysBusMaster_wrData,
  output        sysBusMaster_strb_0,
  output        sysBusMaster_strb_1,
  output        sysBusMaster_strb_2,
  output        sysBusMaster_strb_3
);
  wire [31:0] alu_io_source1; // @[EX.scala 33:19]
  wire [31:0] alu_io_source2; // @[EX.scala 33:19]
  wire [3:0] alu_io_operation; // @[EX.scala 33:19]
  wire [31:0] alu_io_output; // @[EX.scala 33:19]
  wire [2:0] branchControl_io_funct3; // @[EX.scala 34:29]
  wire [31:0] branchControl_io_registerS1; // @[EX.scala 34:29]
  wire [31:0] branchControl_io_registerS2; // @[EX.scala 34:29]
  wire  branchControl_io_jump; // @[EX.scala 34:29]
  wire  branchControl_io_takeBranch; // @[EX.scala 34:29]
  wire [31:0] fwdRegOp1 = ctrl_fwdA_en ? $signed(ctrl_fwdA) : $signed(in_regOp1); // @[EX.scala 35:22]
  wire [31:0] fwdRegOp2 = ctrl_fwdB_en ? $signed(ctrl_fwdB) : $signed(in_regOp2); // @[EX.scala 36:22]
  wire  _T = branchControl_io_takeBranch; // @[EX.scala 43:58]
  wire [31:0] _T_5 = $signed(fwdRegOp1) + $signed(in_imm); // @[EX.scala 44:72]
  wire [31:0] _T_10 = $signed(in_pc) + $signed(in_imm); // @[EX.scala 44:112]
  wire  _T_19 = 2'h0 == in_aluSrc1; // @[Conditional.scala 37:30]
  wire  _T_20 = 2'h1 == in_aluSrc1; // @[Conditional.scala 37:30]
  wire  _T_22 = 2'h2 == in_aluSrc1; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_1 = _T_22 ? $signed(32'sh0) : $signed(fwdRegOp1); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_20 ? $signed(in_pc) : $signed(_GEN_1); // @[Conditional.scala 39:67]
  wire  _T_23 = 2'h0 == in_aluSrc2; // @[Conditional.scala 37:30]
  wire  _T_24 = 2'h1 == in_aluSrc2; // @[Conditional.scala 37:30]
  wire  _T_25 = 2'h2 == in_aluSrc2; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_4 = _T_25 ? $signed(32'sh4) : $signed(fwdRegOp2); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5 = _T_24 ? $signed(in_imm) : $signed(_GEN_4); // @[Conditional.scala 39:67]
  wire  _T_26 = in_mem != 4'h0; // @[EX.scala 80:15]
  wire [31:0] _T_29 = ctrl_fwdB_en ? $signed(ctrl_fwdB) : $signed(in_regOp2); // @[EX.scala 84:46]
  wire  _T_31 = 2'h1 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _T_33 = 2'h2 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _T_35 = 2'h3 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _GEN_11 = _T_33 | _T_35; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_33 ? 1'h0 : _T_35; // @[Conditional.scala 39:67]
  wire  _GEN_15 = _T_31 | _GEN_11; // @[Conditional.scala 40:58]
  wire  _GEN_16 = _T_31 ? 1'h0 : _GEN_11; // @[Conditional.scala 40:58]
  wire  _GEN_17 = _T_31 ? 1'h0 : _GEN_13; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_19 = in_mem[3] ? 2'h2 : 2'h1; // @[EX.scala 82:20]
  wire [31:0] _GEN_20 = in_mem[3] ? _T_29 : 32'h0; // @[EX.scala 82:20]
  wire  _GEN_21 = in_mem[3] & _GEN_15; // @[EX.scala 82:20]
  wire  _GEN_22 = in_mem[3] & _GEN_16; // @[EX.scala 82:20]
  wire  _GEN_23 = in_mem[3] & _GEN_17; // @[EX.scala 82:20]
  ALU alu ( // @[EX.scala 33:19]
    .io_source1(alu_io_source1),
    .io_source2(alu_io_source2),
    .io_operation(alu_io_operation),
    .io_output(alu_io_output)
  );
  BranchControl branchControl ( // @[EX.scala 34:29]
    .io_funct3(branchControl_io_funct3),
    .io_registerS1(branchControl_io_registerS1),
    .io_registerS2(branchControl_io_registerS2),
    .io_jump(branchControl_io_jump),
    .io_takeBranch(branchControl_io_takeBranch)
  );
  assign out_aluRes = alu_io_output; // @[EX.scala 101:14]
  assign out_rd = in_rd; // @[EX.scala 26:10 EX.scala 31:10]
  assign out_wb = in_wb; // @[EX.scala 28:10]
  assign out_wbSrc = in_wbSrc; // @[EX.scala 30:13]
  assign out_mem = in_mem; // @[EX.scala 29:11]
  assign ctrl_rs1 = in_rs1; // @[EX.scala 24:12]
  assign ctrl_rs2 = in_rs2; // @[EX.scala 25:12]
  assign ctrl_rd = in_rd; // @[EX.scala 27:11]
  assign ctrl_branchOut_pcNext = in_brSrc ? _T_5 : _T_10; // @[EX.scala 44:25 EX.scala 48:27]
  assign ctrl_branchOut_branch = _T & in_pcSrc; // @[EX.scala 43:25]
  assign sysBusMaster_cmd = _T_26 ? _GEN_19 : 2'h0; // @[SysBus.scala 57:14 EX.scala 83:24 EX.scala 97:24]
  assign sysBusMaster_addr = _T_26 ? alu_io_output : 32'h0; // @[SysBus.scala 58:15 EX.scala 81:23]
  assign sysBusMaster_wrData = _T_26 ? _GEN_20 : 32'h0; // @[SysBus.scala 59:17 EX.scala 84:27]
  assign sysBusMaster_strb_0 = _T_26 & _GEN_21; // @[SysBus.scala 60:15 EX.scala 87:29 EX.scala 90:29 EX.scala 93:29]
  assign sysBusMaster_strb_1 = _T_26 & _GEN_22; // @[SysBus.scala 60:15 EX.scala 87:29 EX.scala 90:29 EX.scala 93:29]
  assign sysBusMaster_strb_2 = _T_26 & _GEN_23; // @[SysBus.scala 60:15 EX.scala 87:29 EX.scala 90:29 EX.scala 93:29]
  assign sysBusMaster_strb_3 = _T_26 & _GEN_23; // @[SysBus.scala 60:15 EX.scala 87:29 EX.scala 90:29 EX.scala 93:29]
  assign alu_io_source1 = _T_19 ? $signed(fwdRegOp1) : $signed(_GEN_2); // @[EX.scala 51:18 EX.scala 57:22 EX.scala 60:22 EX.scala 63:22]
  assign alu_io_source2 = _T_23 ? $signed(fwdRegOp2) : $signed(_GEN_5); // @[EX.scala 52:18 EX.scala 68:22 EX.scala 71:22 EX.scala 74:22]
  assign alu_io_operation = in_aluOp; // @[EX.scala 53:20]
  assign branchControl_io_funct3 = in_funct3; // @[EX.scala 38:27]
  assign branchControl_io_registerS1 = ctrl_fwdA_en ? $signed(ctrl_fwdA) : $signed(in_regOp1); // @[EX.scala 40:31]
  assign branchControl_io_registerS2 = ctrl_fwdB_en ? $signed(ctrl_fwdB) : $signed(in_regOp2); // @[EX.scala 41:31]
  assign branchControl_io_jump = in_jump; // @[EX.scala 39:25]
endmodule
module MEM(
  input  [31:0] in_aluRes,
  input  [4:0]  in_rd,
  input         in_wb,
  input         in_wbSrc,
  input  [3:0]  in_mem,
  output [31:0] out_memRes,
  output [31:0] out_aluRes,
  output [4:0]  out_rd,
  output        out_wb,
  output        out_wbSrc,
  input  [31:0] sysBusSlave_rdData,
  output [4:0]  ctrl_rd,
  output [31:0] ctrl_aluRes
);
  wire  _T_1 = in_mem != 4'h0; // @[MEM.scala 20:15]
  wire  _T_3 = ~in_mem[3]; // @[MEM.scala 20:26]
  wire  _T_4 = _T_1 & _T_3; // @[MEM.scala 20:23]
  wire [7:0] rdData_0 = _T_4 ? sysBusSlave_rdData[7:0] : 8'h0; // @[MEM.scala 20:37]
  wire [7:0] rdData_1 = _T_4 ? sysBusSlave_rdData[15:8] : 8'h0; // @[MEM.scala 20:37]
  wire [7:0] rdData_2 = _T_4 ? sysBusSlave_rdData[23:16] : 8'h0; // @[MEM.scala 20:37]
  wire [7:0] rdData_3 = _T_4 ? sysBusSlave_rdData[31:24] : 8'h0; // @[MEM.scala 20:37]
  wire  _T_11 = 2'h1 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _T_14 = in_mem[2] & rdData_0[7]; // @[MEM.scala 27:56]
  wire [5:0] _T_89 = {_T_14,_T_14,_T_14,_T_14,_T_14,_T_14}; // @[MEM.scala 27:73]
  wire [11:0] _T_95 = {_T_14,_T_14,_T_14,_T_14,_T_14,_T_14,_T_89}; // @[MEM.scala 27:73]
  wire [31:0] _T_109 = {_T_14,_T_14,_T_14,_T_14,_T_14,_T_14,_T_89,_T_95,rdData_0}; // @[MEM.scala 27:92]
  wire  _T_110 = 2'h2 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire  _T_113 = in_mem[2] & rdData_1[7]; // @[MEM.scala 30:56]
  wire [7:0] _T_166 = {_T_113,_T_113,_T_113,_T_113,_T_113,_T_113,_T_113,_T_113}; // @[MEM.scala 30:73]
  wire [23:0] _T_175 = {_T_113,_T_113,_T_113,_T_113,_T_113,_T_113,_T_113,_T_113,_T_166,rdData_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_177 = {_T_175,rdData_0}; // @[MEM.scala 30:103]
  wire  _T_178 = 2'h3 == in_mem[1:0]; // @[Conditional.scala 37:30]
  wire [31:0] _T_182 = {rdData_3,rdData_2,rdData_1,rdData_0}; // @[MEM.scala 33:72]
  wire [31:0] _GEN_4 = _T_178 ? $signed(_T_182) : $signed(32'sh0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_5 = _T_110 ? $signed(_T_177) : $signed(_GEN_4); // @[Conditional.scala 39:67]
  assign out_memRes = _T_11 ? $signed(_T_109) : $signed(_GEN_5); // @[MEM.scala 24:14 MEM.scala 27:18 MEM.scala 30:18 MEM.scala 33:18]
  assign out_aluRes = in_aluRes; // @[MEM.scala 40:14]
  assign out_rd = in_rd; // @[MEM.scala 39:10]
  assign out_wb = in_wb; // @[MEM.scala 37:10]
  assign out_wbSrc = in_wbSrc; // @[MEM.scala 38:13]
  assign ctrl_rd = in_rd; // @[MEM.scala 42:11]
  assign ctrl_aluRes = in_aluRes; // @[MEM.scala 41:15]
endmodule
module WB(
  input  [31:0] in_memRes,
  input  [31:0] in_aluRes,
  input  [4:0]  in_rd,
  input         in_wb,
  input         in_wbSrc,
  output [4:0]  out_rd,
  output [31:0] out_res,
  output        out_wb,
  output [4:0]  ctrl_rd,
  output [31:0] ctrl_res
);
  assign out_rd = in_rd; // @[WB.scala 17:10]
  assign out_res = in_wbSrc ? $signed(in_memRes) : $signed(in_aluRes); // @[WB.scala 14:11]
  assign out_wb = in_wb; // @[WB.scala 18:10]
  assign ctrl_rd = in_rd; // @[WB.scala 15:11]
  assign ctrl_res = in_wbSrc ? $signed(in_memRes) : $signed(in_aluRes); // @[WB.scala 16:12]
endmodule
module ForwardingUnit(
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd_MEM,
  input         io_wb_MEM,
  input  [4:0]  io_rd_WB,
  input         io_wb_WB,
  input  [31:0] io_aluRes_MEM,
  input  [31:0] io_res_WB,
  output [31:0] io_fwdA,
  output [31:0] io_fwdB,
  output        io_fwdA_en,
  output        io_fwdB_en
);
  wire  _T = io_rs1 == io_rd_MEM; // @[ForwardingUnit.scala 24:15]
  wire  _T_1 = _T & io_wb_MEM; // @[ForwardingUnit.scala 24:29]
  wire  _T_2 = io_rs1 == io_rd_WB; // @[ForwardingUnit.scala 28:21]
  wire  _T_3 = _T_2 & io_wb_WB; // @[ForwardingUnit.scala 28:34]
  wire [31:0] _GEN_1 = _T_3 ? $signed(io_res_WB) : $signed(32'sh0); // @[ForwardingUnit.scala 28:47]
  wire  _T_4 = io_rs2 == io_rd_MEM; // @[ForwardingUnit.scala 36:15]
  wire  _T_5 = _T_4 & io_wb_MEM; // @[ForwardingUnit.scala 36:29]
  wire  _T_6 = io_rs2 == io_rd_WB; // @[ForwardingUnit.scala 40:21]
  wire  _T_7 = _T_6 & io_wb_WB; // @[ForwardingUnit.scala 40:34]
  wire [31:0] _GEN_5 = _T_7 ? $signed(io_res_WB) : $signed(32'sh0); // @[ForwardingUnit.scala 40:47]
  assign io_fwdA = _T_1 ? $signed(io_aluRes_MEM) : $signed(_GEN_1); // @[ForwardingUnit.scala 26:13 ForwardingUnit.scala 30:13 ForwardingUnit.scala 32:13]
  assign io_fwdB = _T_5 ? $signed(io_aluRes_MEM) : $signed(_GEN_5); // @[ForwardingUnit.scala 38:13 ForwardingUnit.scala 42:13 ForwardingUnit.scala 44:13]
  assign io_fwdA_en = _T_1 | _T_3; // @[ForwardingUnit.scala 22:14 ForwardingUnit.scala 25:16 ForwardingUnit.scala 29:16]
  assign io_fwdB_en = _T_5 | _T_7; // @[ForwardingUnit.scala 35:14 ForwardingUnit.scala 37:16 ForwardingUnit.scala 41:16]
endmodule
module HazardDetectionUnit(
  output        io_pcEn,
  output        io_flushIF,
  output        io_flushID,
  output        io_enableIF_ID,
  input  [4:0]  io_rd_EX,
  input  [31:0] io_instr,
  input         io_wbSrc_EX,
  input         io_branch_EX
);
  wire [4:0] rs1 = io_instr[19:15]; // @[HazardDetectionUnit.scala 22:21]
  wire [4:0] rs2 = io_instr[24:20]; // @[HazardDetectionUnit.scala 23:21]
  wire  rs1IsAccessed = io_rd_EX == rs1; // @[HazardDetectionUnit.scala 24:32]
  wire  rs2IsAccessed = io_rd_EX == rs2; // @[HazardDetectionUnit.scala 25:32]
  wire  _T = rs1IsAccessed | rs2IsAccessed; // @[HazardDetectionUnit.scala 26:23]
  wire  _T_1 = _T & io_wbSrc_EX; // @[HazardDetectionUnit.scala 26:41]
  wire  _GEN_0 = _T_1 ? 1'h0 : 1'h1; // @[HazardDetectionUnit.scala 26:57]
  assign io_pcEn = _T_1 ? 1'h0 : 1'h1; // @[HazardDetectionUnit.scala 17:11 HazardDetectionUnit.scala 27:13]
  assign io_flushIF = io_branch_EX; // @[HazardDetectionUnit.scala 18:14 HazardDetectionUnit.scala 33:16]
  assign io_flushID = io_branch_EX | _T_1; // @[HazardDetectionUnit.scala 19:14 HazardDetectionUnit.scala 28:16 HazardDetectionUnit.scala 34:16]
  assign io_enableIF_ID = io_branch_EX ? 1'h0 : _GEN_0; // @[HazardDetectionUnit.scala 20:18 HazardDetectionUnit.scala 29:20 HazardDetectionUnit.scala 35:20]
endmodule
module RVPipeline(
  input         clock,
  input         reset,
  output [1:0]  io_sysBusIO_m_cmd,
  output [31:0] io_sysBusIO_m_addr,
  output [31:0] io_sysBusIO_m_wrData,
  output        io_sysBusIO_m_strb_0,
  output        io_sysBusIO_m_strb_1,
  output        io_sysBusIO_m_strb_2,
  output        io_sysBusIO_m_strb_3,
  input  [31:0] io_sysBusIO_s_rdData,
  output [31:0] io_instrBus_pc,
  input  [31:0] io_instrBus_instr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  ifStage_clock; // @[RVPipeline.scala 18:23]
  wire  ifStage_reset; // @[RVPipeline.scala 18:23]
  wire [31:0] ifStage_in_pcNext; // @[RVPipeline.scala 18:23]
  wire  ifStage_in_branch; // @[RVPipeline.scala 18:23]
  wire [31:0] ifStage_out_pc; // @[RVPipeline.scala 18:23]
  wire [31:0] ifStage_out_instr; // @[RVPipeline.scala 18:23]
  wire [31:0] ifStage_instrBus_pc; // @[RVPipeline.scala 18:23]
  wire [31:0] ifStage_instrBus_instr; // @[RVPipeline.scala 18:23]
  wire  ifStage_ctrl_pcEn; // @[RVPipeline.scala 18:23]
  wire  idStage_clock; // @[RVPipeline.scala 19:23]
  wire  idStage_reset; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_in_pc; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_in_instr; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_out_pc; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_out_imm; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_out_regOp1; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_out_regOp2; // @[RVPipeline.scala 19:23]
  wire [4:0] idStage_out_rs1; // @[RVPipeline.scala 19:23]
  wire [4:0] idStage_out_rs2; // @[RVPipeline.scala 19:23]
  wire [4:0] idStage_out_rd; // @[RVPipeline.scala 19:23]
  wire [3:0] idStage_out_aluOp; // @[RVPipeline.scala 19:23]
  wire [1:0] idStage_out_aluSrc1; // @[RVPipeline.scala 19:23]
  wire [1:0] idStage_out_aluSrc2; // @[RVPipeline.scala 19:23]
  wire  idStage_out_brSrc; // @[RVPipeline.scala 19:23]
  wire  idStage_out_pcSrc; // @[RVPipeline.scala 19:23]
  wire  idStage_out_wb; // @[RVPipeline.scala 19:23]
  wire  idStage_out_wbSrc; // @[RVPipeline.scala 19:23]
  wire [3:0] idStage_out_mem; // @[RVPipeline.scala 19:23]
  wire  idStage_out_jump; // @[RVPipeline.scala 19:23]
  wire [2:0] idStage_out_funct3; // @[RVPipeline.scala 19:23]
  wire [4:0] idStage_wb_rd; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_wb_res; // @[RVPipeline.scala 19:23]
  wire  idStage_wb_wb; // @[RVPipeline.scala 19:23]
  wire  idStage_ctrl_flushID; // @[RVPipeline.scala 19:23]
  wire [31:0] idStage_ctrl_instr; // @[RVPipeline.scala 19:23]
  wire [31:0] exStage_in_pc; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_in_imm; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_in_regOp1; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_in_regOp2; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_in_rs1; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_in_rs2; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_in_rd; // @[RVPipeline.scala 20:23]
  wire [3:0] exStage_in_aluOp; // @[RVPipeline.scala 20:23]
  wire [1:0] exStage_in_aluSrc1; // @[RVPipeline.scala 20:23]
  wire [1:0] exStage_in_aluSrc2; // @[RVPipeline.scala 20:23]
  wire  exStage_in_brSrc; // @[RVPipeline.scala 20:23]
  wire  exStage_in_pcSrc; // @[RVPipeline.scala 20:23]
  wire  exStage_in_wb; // @[RVPipeline.scala 20:23]
  wire  exStage_in_wbSrc; // @[RVPipeline.scala 20:23]
  wire [3:0] exStage_in_mem; // @[RVPipeline.scala 20:23]
  wire  exStage_in_jump; // @[RVPipeline.scala 20:23]
  wire [2:0] exStage_in_funct3; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_out_aluRes; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_out_rd; // @[RVPipeline.scala 20:23]
  wire  exStage_out_wb; // @[RVPipeline.scala 20:23]
  wire  exStage_out_wbSrc; // @[RVPipeline.scala 20:23]
  wire [3:0] exStage_out_mem; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_ctrl_rs1; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_ctrl_rs2; // @[RVPipeline.scala 20:23]
  wire [4:0] exStage_ctrl_rd; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_ctrl_fwdA; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_ctrl_fwdB; // @[RVPipeline.scala 20:23]
  wire  exStage_ctrl_fwdA_en; // @[RVPipeline.scala 20:23]
  wire  exStage_ctrl_fwdB_en; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_ctrl_branchOut_pcNext; // @[RVPipeline.scala 20:23]
  wire  exStage_ctrl_branchOut_branch; // @[RVPipeline.scala 20:23]
  wire [1:0] exStage_sysBusMaster_cmd; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_sysBusMaster_addr; // @[RVPipeline.scala 20:23]
  wire [31:0] exStage_sysBusMaster_wrData; // @[RVPipeline.scala 20:23]
  wire  exStage_sysBusMaster_strb_0; // @[RVPipeline.scala 20:23]
  wire  exStage_sysBusMaster_strb_1; // @[RVPipeline.scala 20:23]
  wire  exStage_sysBusMaster_strb_2; // @[RVPipeline.scala 20:23]
  wire  exStage_sysBusMaster_strb_3; // @[RVPipeline.scala 20:23]
  wire [31:0] memStage_in_aluRes; // @[RVPipeline.scala 21:24]
  wire [4:0] memStage_in_rd; // @[RVPipeline.scala 21:24]
  wire  memStage_in_wb; // @[RVPipeline.scala 21:24]
  wire  memStage_in_wbSrc; // @[RVPipeline.scala 21:24]
  wire [3:0] memStage_in_mem; // @[RVPipeline.scala 21:24]
  wire [31:0] memStage_out_memRes; // @[RVPipeline.scala 21:24]
  wire [31:0] memStage_out_aluRes; // @[RVPipeline.scala 21:24]
  wire [4:0] memStage_out_rd; // @[RVPipeline.scala 21:24]
  wire  memStage_out_wb; // @[RVPipeline.scala 21:24]
  wire  memStage_out_wbSrc; // @[RVPipeline.scala 21:24]
  wire [31:0] memStage_sysBusSlave_rdData; // @[RVPipeline.scala 21:24]
  wire [4:0] memStage_ctrl_rd; // @[RVPipeline.scala 21:24]
  wire [31:0] memStage_ctrl_aluRes; // @[RVPipeline.scala 21:24]
  wire [31:0] wbStage_in_memRes; // @[RVPipeline.scala 22:23]
  wire [31:0] wbStage_in_aluRes; // @[RVPipeline.scala 22:23]
  wire [4:0] wbStage_in_rd; // @[RVPipeline.scala 22:23]
  wire  wbStage_in_wb; // @[RVPipeline.scala 22:23]
  wire  wbStage_in_wbSrc; // @[RVPipeline.scala 22:23]
  wire [4:0] wbStage_out_rd; // @[RVPipeline.scala 22:23]
  wire [31:0] wbStage_out_res; // @[RVPipeline.scala 22:23]
  wire  wbStage_out_wb; // @[RVPipeline.scala 22:23]
  wire [4:0] wbStage_ctrl_rd; // @[RVPipeline.scala 22:23]
  wire [31:0] wbStage_ctrl_res; // @[RVPipeline.scala 22:23]
  wire [4:0] forwardingUnit_io_rs1; // @[RVPipeline.scala 30:30]
  wire [4:0] forwardingUnit_io_rs2; // @[RVPipeline.scala 30:30]
  wire [4:0] forwardingUnit_io_rd_MEM; // @[RVPipeline.scala 30:30]
  wire  forwardingUnit_io_wb_MEM; // @[RVPipeline.scala 30:30]
  wire [4:0] forwardingUnit_io_rd_WB; // @[RVPipeline.scala 30:30]
  wire  forwardingUnit_io_wb_WB; // @[RVPipeline.scala 30:30]
  wire [31:0] forwardingUnit_io_aluRes_MEM; // @[RVPipeline.scala 30:30]
  wire [31:0] forwardingUnit_io_res_WB; // @[RVPipeline.scala 30:30]
  wire [31:0] forwardingUnit_io_fwdA; // @[RVPipeline.scala 30:30]
  wire [31:0] forwardingUnit_io_fwdB; // @[RVPipeline.scala 30:30]
  wire  forwardingUnit_io_fwdA_en; // @[RVPipeline.scala 30:30]
  wire  forwardingUnit_io_fwdB_en; // @[RVPipeline.scala 30:30]
  wire  hazardDetectionUnit_io_pcEn; // @[RVPipeline.scala 31:35]
  wire  hazardDetectionUnit_io_flushIF; // @[RVPipeline.scala 31:35]
  wire  hazardDetectionUnit_io_flushID; // @[RVPipeline.scala 31:35]
  wire  hazardDetectionUnit_io_enableIF_ID; // @[RVPipeline.scala 31:35]
  wire [4:0] hazardDetectionUnit_io_rd_EX; // @[RVPipeline.scala 31:35]
  wire [31:0] hazardDetectionUnit_io_instr; // @[RVPipeline.scala 31:35]
  wire  hazardDetectionUnit_io_wbSrc_EX; // @[RVPipeline.scala 31:35]
  wire  hazardDetectionUnit_io_branch_EX; // @[RVPipeline.scala 31:35]
  reg [31:0] if_id_pc; // @[RVPipeline.scala 33:22]
  reg [31:0] if_id_instr; // @[RVPipeline.scala 33:22]
  reg [31:0] id_ex_pc; // @[RVPipeline.scala 34:22]
  reg [31:0] id_ex_imm; // @[RVPipeline.scala 34:22]
  reg [31:0] id_ex_regOp1; // @[RVPipeline.scala 34:22]
  reg [31:0] id_ex_regOp2; // @[RVPipeline.scala 34:22]
  reg [4:0] id_ex_rs1; // @[RVPipeline.scala 34:22]
  reg [4:0] id_ex_rs2; // @[RVPipeline.scala 34:22]
  reg [4:0] id_ex_rd; // @[RVPipeline.scala 34:22]
  reg [3:0] id_ex_aluOp; // @[RVPipeline.scala 34:22]
  reg [1:0] id_ex_aluSrc1; // @[RVPipeline.scala 34:22]
  reg [1:0] id_ex_aluSrc2; // @[RVPipeline.scala 34:22]
  reg  id_ex_brSrc; // @[RVPipeline.scala 34:22]
  reg  id_ex_pcSrc; // @[RVPipeline.scala 34:22]
  reg  id_ex_wb; // @[RVPipeline.scala 34:22]
  reg  id_ex_wbSrc; // @[RVPipeline.scala 34:22]
  reg [3:0] id_ex_mem; // @[RVPipeline.scala 34:22]
  reg  id_ex_jump; // @[RVPipeline.scala 34:22]
  reg [2:0] id_ex_funct3; // @[RVPipeline.scala 34:22]
  reg [31:0] ex_mem_aluRes; // @[RVPipeline.scala 35:23]
  reg [4:0] ex_mem_rd; // @[RVPipeline.scala 35:23]
  reg  ex_mem_wb; // @[RVPipeline.scala 35:23]
  reg  ex_mem_wbSrc; // @[RVPipeline.scala 35:23]
  reg [3:0] ex_mem_mem; // @[RVPipeline.scala 35:23]
  reg [31:0] mem_wb_memRes; // @[RVPipeline.scala 36:23]
  reg [31:0] mem_wb_aluRes; // @[RVPipeline.scala 36:23]
  reg [4:0] mem_wb_rd; // @[RVPipeline.scala 36:23]
  reg  mem_wb_wb; // @[RVPipeline.scala 36:23]
  reg  mem_wb_wbSrc; // @[RVPipeline.scala 36:23]
  IF ifStage ( // @[RVPipeline.scala 18:23]
    .clock(ifStage_clock),
    .reset(ifStage_reset),
    .in_pcNext(ifStage_in_pcNext),
    .in_branch(ifStage_in_branch),
    .out_pc(ifStage_out_pc),
    .out_instr(ifStage_out_instr),
    .instrBus_pc(ifStage_instrBus_pc),
    .instrBus_instr(ifStage_instrBus_instr),
    .ctrl_pcEn(ifStage_ctrl_pcEn)
  );
  ID idStage ( // @[RVPipeline.scala 19:23]
    .clock(idStage_clock),
    .reset(idStage_reset),
    .in_pc(idStage_in_pc),
    .in_instr(idStage_in_instr),
    .out_pc(idStage_out_pc),
    .out_imm(idStage_out_imm),
    .out_regOp1(idStage_out_regOp1),
    .out_regOp2(idStage_out_regOp2),
    .out_rs1(idStage_out_rs1),
    .out_rs2(idStage_out_rs2),
    .out_rd(idStage_out_rd),
    .out_aluOp(idStage_out_aluOp),
    .out_aluSrc1(idStage_out_aluSrc1),
    .out_aluSrc2(idStage_out_aluSrc2),
    .out_brSrc(idStage_out_brSrc),
    .out_pcSrc(idStage_out_pcSrc),
    .out_wb(idStage_out_wb),
    .out_wbSrc(idStage_out_wbSrc),
    .out_mem(idStage_out_mem),
    .out_jump(idStage_out_jump),
    .out_funct3(idStage_out_funct3),
    .wb_rd(idStage_wb_rd),
    .wb_res(idStage_wb_res),
    .wb_wb(idStage_wb_wb),
    .ctrl_flushID(idStage_ctrl_flushID),
    .ctrl_instr(idStage_ctrl_instr)
  );
  EX exStage ( // @[RVPipeline.scala 20:23]
    .in_pc(exStage_in_pc),
    .in_imm(exStage_in_imm),
    .in_regOp1(exStage_in_regOp1),
    .in_regOp2(exStage_in_regOp2),
    .in_rs1(exStage_in_rs1),
    .in_rs2(exStage_in_rs2),
    .in_rd(exStage_in_rd),
    .in_aluOp(exStage_in_aluOp),
    .in_aluSrc1(exStage_in_aluSrc1),
    .in_aluSrc2(exStage_in_aluSrc2),
    .in_brSrc(exStage_in_brSrc),
    .in_pcSrc(exStage_in_pcSrc),
    .in_wb(exStage_in_wb),
    .in_wbSrc(exStage_in_wbSrc),
    .in_mem(exStage_in_mem),
    .in_jump(exStage_in_jump),
    .in_funct3(exStage_in_funct3),
    .out_aluRes(exStage_out_aluRes),
    .out_rd(exStage_out_rd),
    .out_wb(exStage_out_wb),
    .out_wbSrc(exStage_out_wbSrc),
    .out_mem(exStage_out_mem),
    .ctrl_rs1(exStage_ctrl_rs1),
    .ctrl_rs2(exStage_ctrl_rs2),
    .ctrl_rd(exStage_ctrl_rd),
    .ctrl_fwdA(exStage_ctrl_fwdA),
    .ctrl_fwdB(exStage_ctrl_fwdB),
    .ctrl_fwdA_en(exStage_ctrl_fwdA_en),
    .ctrl_fwdB_en(exStage_ctrl_fwdB_en),
    .ctrl_branchOut_pcNext(exStage_ctrl_branchOut_pcNext),
    .ctrl_branchOut_branch(exStage_ctrl_branchOut_branch),
    .sysBusMaster_cmd(exStage_sysBusMaster_cmd),
    .sysBusMaster_addr(exStage_sysBusMaster_addr),
    .sysBusMaster_wrData(exStage_sysBusMaster_wrData),
    .sysBusMaster_strb_0(exStage_sysBusMaster_strb_0),
    .sysBusMaster_strb_1(exStage_sysBusMaster_strb_1),
    .sysBusMaster_strb_2(exStage_sysBusMaster_strb_2),
    .sysBusMaster_strb_3(exStage_sysBusMaster_strb_3)
  );
  MEM memStage ( // @[RVPipeline.scala 21:24]
    .in_aluRes(memStage_in_aluRes),
    .in_rd(memStage_in_rd),
    .in_wb(memStage_in_wb),
    .in_wbSrc(memStage_in_wbSrc),
    .in_mem(memStage_in_mem),
    .out_memRes(memStage_out_memRes),
    .out_aluRes(memStage_out_aluRes),
    .out_rd(memStage_out_rd),
    .out_wb(memStage_out_wb),
    .out_wbSrc(memStage_out_wbSrc),
    .sysBusSlave_rdData(memStage_sysBusSlave_rdData),
    .ctrl_rd(memStage_ctrl_rd),
    .ctrl_aluRes(memStage_ctrl_aluRes)
  );
  WB wbStage ( // @[RVPipeline.scala 22:23]
    .in_memRes(wbStage_in_memRes),
    .in_aluRes(wbStage_in_aluRes),
    .in_rd(wbStage_in_rd),
    .in_wb(wbStage_in_wb),
    .in_wbSrc(wbStage_in_wbSrc),
    .out_rd(wbStage_out_rd),
    .out_res(wbStage_out_res),
    .out_wb(wbStage_out_wb),
    .ctrl_rd(wbStage_ctrl_rd),
    .ctrl_res(wbStage_ctrl_res)
  );
  ForwardingUnit forwardingUnit ( // @[RVPipeline.scala 30:30]
    .io_rs1(forwardingUnit_io_rs1),
    .io_rs2(forwardingUnit_io_rs2),
    .io_rd_MEM(forwardingUnit_io_rd_MEM),
    .io_wb_MEM(forwardingUnit_io_wb_MEM),
    .io_rd_WB(forwardingUnit_io_rd_WB),
    .io_wb_WB(forwardingUnit_io_wb_WB),
    .io_aluRes_MEM(forwardingUnit_io_aluRes_MEM),
    .io_res_WB(forwardingUnit_io_res_WB),
    .io_fwdA(forwardingUnit_io_fwdA),
    .io_fwdB(forwardingUnit_io_fwdB),
    .io_fwdA_en(forwardingUnit_io_fwdA_en),
    .io_fwdB_en(forwardingUnit_io_fwdB_en)
  );
  HazardDetectionUnit hazardDetectionUnit ( // @[RVPipeline.scala 31:35]
    .io_pcEn(hazardDetectionUnit_io_pcEn),
    .io_flushIF(hazardDetectionUnit_io_flushIF),
    .io_flushID(hazardDetectionUnit_io_flushID),
    .io_enableIF_ID(hazardDetectionUnit_io_enableIF_ID),
    .io_rd_EX(hazardDetectionUnit_io_rd_EX),
    .io_instr(hazardDetectionUnit_io_instr),
    .io_wbSrc_EX(hazardDetectionUnit_io_wbSrc_EX),
    .io_branch_EX(hazardDetectionUnit_io_branch_EX)
  );
  assign io_sysBusIO_m_cmd = exStage_sysBusMaster_cmd; // @[RVPipeline.scala 81:17]
  assign io_sysBusIO_m_addr = exStage_sysBusMaster_addr; // @[RVPipeline.scala 81:17]
  assign io_sysBusIO_m_wrData = exStage_sysBusMaster_wrData; // @[RVPipeline.scala 81:17]
  assign io_sysBusIO_m_strb_0 = exStage_sysBusMaster_strb_0; // @[RVPipeline.scala 81:17]
  assign io_sysBusIO_m_strb_1 = exStage_sysBusMaster_strb_1; // @[RVPipeline.scala 81:17]
  assign io_sysBusIO_m_strb_2 = exStage_sysBusMaster_strb_2; // @[RVPipeline.scala 81:17]
  assign io_sysBusIO_m_strb_3 = exStage_sysBusMaster_strb_3; // @[RVPipeline.scala 81:17]
  assign io_instrBus_pc = ifStage_instrBus_pc; // @[RVPipeline.scala 39:20]
  assign ifStage_clock = clock;
  assign ifStage_reset = reset;
  assign ifStage_in_pcNext = exStage_ctrl_branchOut_pcNext; // @[RVPipeline.scala 40:14]
  assign ifStage_in_branch = exStage_ctrl_branchOut_branch; // @[RVPipeline.scala 40:14]
  assign ifStage_instrBus_instr = io_instrBus_instr; // @[RVPipeline.scala 39:20]
  assign ifStage_ctrl_pcEn = hazardDetectionUnit_io_pcEn; // @[RVPipeline.scala 41:21]
  assign idStage_clock = clock;
  assign idStage_reset = reset;
  assign idStage_in_pc = if_id_pc; // @[RVPipeline.scala 50:14]
  assign idStage_in_instr = if_id_instr; // @[RVPipeline.scala 50:14]
  assign idStage_wb_rd = wbStage_out_rd; // @[RVPipeline.scala 49:14]
  assign idStage_wb_res = wbStage_out_res; // @[RVPipeline.scala 49:14]
  assign idStage_wb_wb = wbStage_out_wb; // @[RVPipeline.scala 49:14]
  assign idStage_ctrl_flushID = hazardDetectionUnit_io_flushID; // @[RVPipeline.scala 48:24]
  assign exStage_in_pc = id_ex_pc; // @[RVPipeline.scala 55:14]
  assign exStage_in_imm = id_ex_imm; // @[RVPipeline.scala 55:14]
  assign exStage_in_regOp1 = id_ex_regOp1; // @[RVPipeline.scala 55:14]
  assign exStage_in_regOp2 = id_ex_regOp2; // @[RVPipeline.scala 55:14]
  assign exStage_in_rs1 = id_ex_rs1; // @[RVPipeline.scala 55:14]
  assign exStage_in_rs2 = id_ex_rs2; // @[RVPipeline.scala 55:14]
  assign exStage_in_rd = id_ex_rd; // @[RVPipeline.scala 55:14]
  assign exStage_in_aluOp = id_ex_aluOp; // @[RVPipeline.scala 55:14]
  assign exStage_in_aluSrc1 = id_ex_aluSrc1; // @[RVPipeline.scala 55:14]
  assign exStage_in_aluSrc2 = id_ex_aluSrc2; // @[RVPipeline.scala 55:14]
  assign exStage_in_brSrc = id_ex_brSrc; // @[RVPipeline.scala 55:14]
  assign exStage_in_pcSrc = id_ex_pcSrc; // @[RVPipeline.scala 55:14]
  assign exStage_in_wb = id_ex_wb; // @[RVPipeline.scala 55:14]
  assign exStage_in_wbSrc = id_ex_wbSrc; // @[RVPipeline.scala 55:14]
  assign exStage_in_mem = id_ex_mem; // @[RVPipeline.scala 55:14]
  assign exStage_in_jump = id_ex_jump; // @[RVPipeline.scala 55:14]
  assign exStage_in_funct3 = id_ex_funct3; // @[RVPipeline.scala 55:14]
  assign exStage_ctrl_fwdA = forwardingUnit_io_fwdA; // @[RVPipeline.scala 62:21]
  assign exStage_ctrl_fwdB = forwardingUnit_io_fwdB; // @[RVPipeline.scala 63:21]
  assign exStage_ctrl_fwdA_en = forwardingUnit_io_fwdA_en; // @[RVPipeline.scala 64:24]
  assign exStage_ctrl_fwdB_en = forwardingUnit_io_fwdB_en; // @[RVPipeline.scala 65:24]
  assign memStage_in_aluRes = ex_mem_aluRes; // @[RVPipeline.scala 69:15]
  assign memStage_in_rd = ex_mem_rd; // @[RVPipeline.scala 69:15]
  assign memStage_in_wb = ex_mem_wb; // @[RVPipeline.scala 69:15]
  assign memStage_in_wbSrc = ex_mem_wbSrc; // @[RVPipeline.scala 69:15]
  assign memStage_in_mem = ex_mem_mem; // @[RVPipeline.scala 69:15]
  assign memStage_sysBusSlave_rdData = io_sysBusIO_s_rdData; // @[RVPipeline.scala 82:17]
  assign wbStage_in_memRes = mem_wb_memRes; // @[RVPipeline.scala 76:14]
  assign wbStage_in_aluRes = mem_wb_aluRes; // @[RVPipeline.scala 76:14]
  assign wbStage_in_rd = mem_wb_rd; // @[RVPipeline.scala 76:14]
  assign wbStage_in_wb = mem_wb_wb; // @[RVPipeline.scala 76:14]
  assign wbStage_in_wbSrc = mem_wb_wbSrc; // @[RVPipeline.scala 76:14]
  assign forwardingUnit_io_rs1 = exStage_ctrl_rs1; // @[RVPipeline.scala 57:25]
  assign forwardingUnit_io_rs2 = exStage_ctrl_rs2; // @[RVPipeline.scala 58:25]
  assign forwardingUnit_io_rd_MEM = memStage_ctrl_rd; // @[RVPipeline.scala 71:28]
  assign forwardingUnit_io_wb_MEM = memStage_out_wb; // @[RVPipeline.scala 73:28]
  assign forwardingUnit_io_rd_WB = wbStage_ctrl_rd; // @[RVPipeline.scala 77:27]
  assign forwardingUnit_io_wb_WB = wbStage_out_wb; // @[RVPipeline.scala 79:27]
  assign forwardingUnit_io_aluRes_MEM = memStage_ctrl_aluRes; // @[RVPipeline.scala 72:32]
  assign forwardingUnit_io_res_WB = wbStage_ctrl_res; // @[RVPipeline.scala 78:28]
  assign hazardDetectionUnit_io_rd_EX = exStage_ctrl_rd; // @[RVPipeline.scala 59:32]
  assign hazardDetectionUnit_io_instr = idStage_ctrl_instr; // @[RVPipeline.scala 47:32]
  assign hazardDetectionUnit_io_wbSrc_EX = exStage_out_wbSrc; // @[RVPipeline.scala 61:35]
  assign hazardDetectionUnit_io_branch_EX = exStage_ctrl_branchOut_branch; // @[RVPipeline.scala 60:36]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_id_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  if_id_instr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  id_ex_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  id_ex_imm = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  id_ex_regOp1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  id_ex_regOp2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  id_ex_rs1 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  id_ex_rs2 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  id_ex_rd = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  id_ex_aluOp = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  id_ex_aluSrc1 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  id_ex_aluSrc2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  id_ex_brSrc = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  id_ex_pcSrc = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  id_ex_wb = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  id_ex_wbSrc = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  id_ex_mem = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  id_ex_jump = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  id_ex_funct3 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  ex_mem_aluRes = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  ex_mem_rd = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  ex_mem_wb = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ex_mem_wbSrc = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ex_mem_mem = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  mem_wb_memRes = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_wb_aluRes = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_wb_rd = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  mem_wb_wb = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mem_wb_wbSrc = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      if_id_pc <= 32'h0;
    end else if (hazardDetectionUnit_io_flushIF) begin
      if_id_pc <= 32'h0;
    end else if (hazardDetectionUnit_io_enableIF_ID) begin
      if_id_pc <= ifStage_out_pc;
    end
    if (reset) begin
      if_id_instr <= 32'sh0;
    end else if (hazardDetectionUnit_io_flushIF) begin
      if_id_instr <= 32'sh0;
    end else if (hazardDetectionUnit_io_enableIF_ID) begin
      if_id_instr <= ifStage_out_instr;
    end
    if (reset) begin
      id_ex_pc <= 32'h0;
    end else begin
      id_ex_pc <= idStage_out_pc;
    end
    if (reset) begin
      id_ex_imm <= 32'sh0;
    end else begin
      id_ex_imm <= idStage_out_imm;
    end
    if (reset) begin
      id_ex_regOp1 <= 32'sh0;
    end else begin
      id_ex_regOp1 <= idStage_out_regOp1;
    end
    if (reset) begin
      id_ex_regOp2 <= 32'sh0;
    end else begin
      id_ex_regOp2 <= idStage_out_regOp2;
    end
    if (reset) begin
      id_ex_rs1 <= 5'h0;
    end else begin
      id_ex_rs1 <= idStage_out_rs1;
    end
    if (reset) begin
      id_ex_rs2 <= 5'h0;
    end else begin
      id_ex_rs2 <= idStage_out_rs2;
    end
    if (reset) begin
      id_ex_rd <= 5'h0;
    end else begin
      id_ex_rd <= idStage_out_rd;
    end
    if (reset) begin
      id_ex_aluOp <= 4'h0;
    end else begin
      id_ex_aluOp <= idStage_out_aluOp;
    end
    if (reset) begin
      id_ex_aluSrc1 <= 2'h0;
    end else begin
      id_ex_aluSrc1 <= idStage_out_aluSrc1;
    end
    if (reset) begin
      id_ex_aluSrc2 <= 2'h0;
    end else begin
      id_ex_aluSrc2 <= idStage_out_aluSrc2;
    end
    if (reset) begin
      id_ex_brSrc <= 1'h0;
    end else begin
      id_ex_brSrc <= idStage_out_brSrc;
    end
    if (reset) begin
      id_ex_pcSrc <= 1'h0;
    end else begin
      id_ex_pcSrc <= idStage_out_pcSrc;
    end
    if (reset) begin
      id_ex_wb <= 1'h0;
    end else begin
      id_ex_wb <= idStage_out_wb;
    end
    if (reset) begin
      id_ex_wbSrc <= 1'h0;
    end else begin
      id_ex_wbSrc <= idStage_out_wbSrc;
    end
    if (reset) begin
      id_ex_mem <= 4'h0;
    end else begin
      id_ex_mem <= idStage_out_mem;
    end
    if (reset) begin
      id_ex_jump <= 1'h0;
    end else begin
      id_ex_jump <= idStage_out_jump;
    end
    if (reset) begin
      id_ex_funct3 <= 3'h0;
    end else begin
      id_ex_funct3 <= idStage_out_funct3;
    end
    if (reset) begin
      ex_mem_aluRes <= 32'sh0;
    end else begin
      ex_mem_aluRes <= exStage_out_aluRes;
    end
    if (reset) begin
      ex_mem_rd <= 5'h0;
    end else begin
      ex_mem_rd <= exStage_out_rd;
    end
    if (reset) begin
      ex_mem_wb <= 1'h0;
    end else begin
      ex_mem_wb <= exStage_out_wb;
    end
    if (reset) begin
      ex_mem_wbSrc <= 1'h0;
    end else begin
      ex_mem_wbSrc <= exStage_out_wbSrc;
    end
    if (reset) begin
      ex_mem_mem <= 4'h0;
    end else begin
      ex_mem_mem <= exStage_out_mem;
    end
    if (reset) begin
      mem_wb_memRes <= 32'sh0;
    end else begin
      mem_wb_memRes <= memStage_out_memRes;
    end
    if (reset) begin
      mem_wb_aluRes <= 32'sh0;
    end else begin
      mem_wb_aluRes <= memStage_out_aluRes;
    end
    if (reset) begin
      mem_wb_rd <= 5'h0;
    end else begin
      mem_wb_rd <= memStage_out_rd;
    end
    if (reset) begin
      mem_wb_wb <= 1'h0;
    end else begin
      mem_wb_wb <= memStage_out_wb;
    end
    if (reset) begin
      mem_wb_wbSrc <= 1'h0;
    end else begin
      mem_wb_wbSrc <= memStage_out_wbSrc;
    end
  end
endmodule
module ROM(
  input         clock,
  input  [1:0]  sysBusIO_m_cmd,
  input  [31:0] sysBusIO_m_addr,
  output [31:0] sysBusIO_s_rdData,
  input  [31:0] instrBus_pc,
  output [31:0] instrBus_instr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _T_1 = instrBus_pc + 32'h3; // @[ROM.scala 24:42]
  wire [31:0] _T_4 = instrBus_pc + 32'h2; // @[ROM.scala 24:67]
  wire [31:0] _T_7 = instrBus_pc + 32'h1; // @[ROM.scala 24:92]
  wire [7:0] _GEN_1 = 8'h1 == _T_7[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_2 = 8'h2 == _T_7[7:0] ? 8'h0 : _GEN_1; // @[Cat.scala 29:58]
  wire [7:0] _GEN_3 = 8'h3 == _T_7[7:0] ? 8'hfe : _GEN_2; // @[Cat.scala 29:58]
  wire [7:0] _GEN_4 = 8'h4 == _T_7[7:0] ? 8'h93 : _GEN_3; // @[Cat.scala 29:58]
  wire [7:0] _GEN_5 = 8'h5 == _T_7[7:0] ? 8'h5 : _GEN_4; // @[Cat.scala 29:58]
  wire [7:0] _GEN_6 = 8'h6 == _T_7[7:0] ? 8'h0 : _GEN_5; // @[Cat.scala 29:58]
  wire [7:0] _GEN_7 = 8'h7 == _T_7[7:0] ? 8'hfc : _GEN_6; // @[Cat.scala 29:58]
  wire [7:0] _GEN_8 = 8'h8 == _T_7[7:0] ? 8'h33 : _GEN_7; // @[Cat.scala 29:58]
  wire [7:0] _GEN_9 = 8'h9 == _T_7[7:0] ? 8'h6 : _GEN_8; // @[Cat.scala 29:58]
  wire [7:0] _GEN_10 = 8'ha == _T_7[7:0] ? 8'hb5 : _GEN_9; // @[Cat.scala 29:58]
  wire [7:0] _GEN_11 = 8'hb == _T_7[7:0] ? 8'h0 : _GEN_10; // @[Cat.scala 29:58]
  wire [7:0] _GEN_12 = 8'hc == _T_7[7:0] ? 8'h13 : _GEN_11; // @[Cat.scala 29:58]
  wire [7:0] _GEN_13 = 8'hd == _T_7[7:0] ? 8'h5 : _GEN_12; // @[Cat.scala 29:58]
  wire [7:0] _GEN_14 = 8'he == _T_7[7:0] ? 8'ha0 : _GEN_13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_15 = 8'hf == _T_7[7:0] ? 8'h0 : _GEN_14; // @[Cat.scala 29:58]
  wire [7:0] _GEN_16 = 8'h10 == _T_7[7:0] ? 8'h73 : _GEN_15; // @[Cat.scala 29:58]
  wire [7:0] _GEN_17 = 8'h11 == _T_7[7:0] ? 8'h0 : _GEN_16; // @[Cat.scala 29:58]
  wire [7:0] _GEN_18 = 8'h12 == _T_7[7:0] ? 8'h0 : _GEN_17; // @[Cat.scala 29:58]
  wire [7:0] _GEN_19 = 8'h13 == _T_7[7:0] ? 8'h0 : _GEN_18; // @[Cat.scala 29:58]
  wire [7:0] _GEN_20 = 8'h14 == _T_7[7:0] ? 8'h0 : _GEN_19; // @[Cat.scala 29:58]
  wire [7:0] _GEN_21 = 8'h15 == _T_7[7:0] ? 8'h0 : _GEN_20; // @[Cat.scala 29:58]
  wire [7:0] _GEN_22 = 8'h16 == _T_7[7:0] ? 8'h0 : _GEN_21; // @[Cat.scala 29:58]
  wire [7:0] _GEN_23 = 8'h17 == _T_7[7:0] ? 8'h0 : _GEN_22; // @[Cat.scala 29:58]
  wire [7:0] _GEN_24 = 8'h18 == _T_7[7:0] ? 8'h0 : _GEN_23; // @[Cat.scala 29:58]
  wire [7:0] _GEN_25 = 8'h19 == _T_7[7:0] ? 8'h0 : _GEN_24; // @[Cat.scala 29:58]
  wire [7:0] _GEN_26 = 8'h1a == _T_7[7:0] ? 8'h0 : _GEN_25; // @[Cat.scala 29:58]
  wire [7:0] _GEN_27 = 8'h1b == _T_7[7:0] ? 8'h0 : _GEN_26; // @[Cat.scala 29:58]
  wire [7:0] _GEN_28 = 8'h1c == _T_7[7:0] ? 8'h0 : _GEN_27; // @[Cat.scala 29:58]
  wire [7:0] _GEN_29 = 8'h1d == _T_7[7:0] ? 8'h0 : _GEN_28; // @[Cat.scala 29:58]
  wire [7:0] _GEN_30 = 8'h1e == _T_7[7:0] ? 8'h0 : _GEN_29; // @[Cat.scala 29:58]
  wire [7:0] _GEN_31 = 8'h1f == _T_7[7:0] ? 8'h0 : _GEN_30; // @[Cat.scala 29:58]
  wire [7:0] _GEN_32 = 8'h20 == _T_7[7:0] ? 8'h0 : _GEN_31; // @[Cat.scala 29:58]
  wire [7:0] _GEN_33 = 8'h21 == _T_7[7:0] ? 8'h0 : _GEN_32; // @[Cat.scala 29:58]
  wire [7:0] _GEN_34 = 8'h22 == _T_7[7:0] ? 8'h0 : _GEN_33; // @[Cat.scala 29:58]
  wire [7:0] _GEN_35 = 8'h23 == _T_7[7:0] ? 8'h0 : _GEN_34; // @[Cat.scala 29:58]
  wire [7:0] _GEN_36 = 8'h24 == _T_7[7:0] ? 8'h0 : _GEN_35; // @[Cat.scala 29:58]
  wire [7:0] _GEN_37 = 8'h25 == _T_7[7:0] ? 8'h0 : _GEN_36; // @[Cat.scala 29:58]
  wire [7:0] _GEN_38 = 8'h26 == _T_7[7:0] ? 8'h0 : _GEN_37; // @[Cat.scala 29:58]
  wire [7:0] _GEN_39 = 8'h27 == _T_7[7:0] ? 8'h0 : _GEN_38; // @[Cat.scala 29:58]
  wire [7:0] _GEN_40 = 8'h28 == _T_7[7:0] ? 8'h0 : _GEN_39; // @[Cat.scala 29:58]
  wire [7:0] _GEN_41 = 8'h29 == _T_7[7:0] ? 8'h0 : _GEN_40; // @[Cat.scala 29:58]
  wire [7:0] _GEN_42 = 8'h2a == _T_7[7:0] ? 8'h0 : _GEN_41; // @[Cat.scala 29:58]
  wire [7:0] _GEN_43 = 8'h2b == _T_7[7:0] ? 8'h0 : _GEN_42; // @[Cat.scala 29:58]
  wire [7:0] _GEN_44 = 8'h2c == _T_7[7:0] ? 8'h0 : _GEN_43; // @[Cat.scala 29:58]
  wire [7:0] _GEN_45 = 8'h2d == _T_7[7:0] ? 8'h0 : _GEN_44; // @[Cat.scala 29:58]
  wire [7:0] _GEN_46 = 8'h2e == _T_7[7:0] ? 8'h0 : _GEN_45; // @[Cat.scala 29:58]
  wire [7:0] _GEN_47 = 8'h2f == _T_7[7:0] ? 8'h0 : _GEN_46; // @[Cat.scala 29:58]
  wire [7:0] _GEN_48 = 8'h30 == _T_7[7:0] ? 8'h0 : _GEN_47; // @[Cat.scala 29:58]
  wire [7:0] _GEN_49 = 8'h31 == _T_7[7:0] ? 8'h0 : _GEN_48; // @[Cat.scala 29:58]
  wire [7:0] _GEN_50 = 8'h32 == _T_7[7:0] ? 8'h0 : _GEN_49; // @[Cat.scala 29:58]
  wire [7:0] _GEN_51 = 8'h33 == _T_7[7:0] ? 8'h0 : _GEN_50; // @[Cat.scala 29:58]
  wire [7:0] _GEN_52 = 8'h34 == _T_7[7:0] ? 8'h0 : _GEN_51; // @[Cat.scala 29:58]
  wire [7:0] _GEN_53 = 8'h35 == _T_7[7:0] ? 8'h0 : _GEN_52; // @[Cat.scala 29:58]
  wire [7:0] _GEN_54 = 8'h36 == _T_7[7:0] ? 8'h0 : _GEN_53; // @[Cat.scala 29:58]
  wire [7:0] _GEN_55 = 8'h37 == _T_7[7:0] ? 8'h0 : _GEN_54; // @[Cat.scala 29:58]
  wire [7:0] _GEN_56 = 8'h38 == _T_7[7:0] ? 8'h0 : _GEN_55; // @[Cat.scala 29:58]
  wire [7:0] _GEN_57 = 8'h39 == _T_7[7:0] ? 8'h0 : _GEN_56; // @[Cat.scala 29:58]
  wire [7:0] _GEN_58 = 8'h3a == _T_7[7:0] ? 8'h0 : _GEN_57; // @[Cat.scala 29:58]
  wire [7:0] _GEN_59 = 8'h3b == _T_7[7:0] ? 8'h0 : _GEN_58; // @[Cat.scala 29:58]
  wire [7:0] _GEN_60 = 8'h3c == _T_7[7:0] ? 8'h0 : _GEN_59; // @[Cat.scala 29:58]
  wire [7:0] _GEN_61 = 8'h3d == _T_7[7:0] ? 8'h0 : _GEN_60; // @[Cat.scala 29:58]
  wire [7:0] _GEN_62 = 8'h3e == _T_7[7:0] ? 8'h0 : _GEN_61; // @[Cat.scala 29:58]
  wire [7:0] _GEN_63 = 8'h3f == _T_7[7:0] ? 8'h0 : _GEN_62; // @[Cat.scala 29:58]
  wire [7:0] _GEN_64 = 8'h40 == _T_7[7:0] ? 8'h0 : _GEN_63; // @[Cat.scala 29:58]
  wire [7:0] _GEN_65 = 8'h41 == _T_7[7:0] ? 8'h0 : _GEN_64; // @[Cat.scala 29:58]
  wire [7:0] _GEN_66 = 8'h42 == _T_7[7:0] ? 8'h0 : _GEN_65; // @[Cat.scala 29:58]
  wire [7:0] _GEN_67 = 8'h43 == _T_7[7:0] ? 8'h0 : _GEN_66; // @[Cat.scala 29:58]
  wire [7:0] _GEN_68 = 8'h44 == _T_7[7:0] ? 8'h0 : _GEN_67; // @[Cat.scala 29:58]
  wire [7:0] _GEN_69 = 8'h45 == _T_7[7:0] ? 8'h0 : _GEN_68; // @[Cat.scala 29:58]
  wire [7:0] _GEN_70 = 8'h46 == _T_7[7:0] ? 8'h0 : _GEN_69; // @[Cat.scala 29:58]
  wire [7:0] _GEN_71 = 8'h47 == _T_7[7:0] ? 8'h0 : _GEN_70; // @[Cat.scala 29:58]
  wire [7:0] _GEN_72 = 8'h48 == _T_7[7:0] ? 8'h0 : _GEN_71; // @[Cat.scala 29:58]
  wire [7:0] _GEN_73 = 8'h49 == _T_7[7:0] ? 8'h0 : _GEN_72; // @[Cat.scala 29:58]
  wire [7:0] _GEN_74 = 8'h4a == _T_7[7:0] ? 8'h0 : _GEN_73; // @[Cat.scala 29:58]
  wire [7:0] _GEN_75 = 8'h4b == _T_7[7:0] ? 8'h0 : _GEN_74; // @[Cat.scala 29:58]
  wire [7:0] _GEN_76 = 8'h4c == _T_7[7:0] ? 8'h0 : _GEN_75; // @[Cat.scala 29:58]
  wire [7:0] _GEN_77 = 8'h4d == _T_7[7:0] ? 8'h0 : _GEN_76; // @[Cat.scala 29:58]
  wire [7:0] _GEN_78 = 8'h4e == _T_7[7:0] ? 8'h0 : _GEN_77; // @[Cat.scala 29:58]
  wire [7:0] _GEN_79 = 8'h4f == _T_7[7:0] ? 8'h0 : _GEN_78; // @[Cat.scala 29:58]
  wire [7:0] _GEN_80 = 8'h50 == _T_7[7:0] ? 8'h0 : _GEN_79; // @[Cat.scala 29:58]
  wire [7:0] _GEN_81 = 8'h51 == _T_7[7:0] ? 8'h0 : _GEN_80; // @[Cat.scala 29:58]
  wire [7:0] _GEN_82 = 8'h52 == _T_7[7:0] ? 8'h0 : _GEN_81; // @[Cat.scala 29:58]
  wire [7:0] _GEN_83 = 8'h53 == _T_7[7:0] ? 8'h0 : _GEN_82; // @[Cat.scala 29:58]
  wire [7:0] _GEN_84 = 8'h54 == _T_7[7:0] ? 8'h0 : _GEN_83; // @[Cat.scala 29:58]
  wire [7:0] _GEN_85 = 8'h55 == _T_7[7:0] ? 8'h0 : _GEN_84; // @[Cat.scala 29:58]
  wire [7:0] _GEN_86 = 8'h56 == _T_7[7:0] ? 8'h0 : _GEN_85; // @[Cat.scala 29:58]
  wire [7:0] _GEN_87 = 8'h57 == _T_7[7:0] ? 8'h0 : _GEN_86; // @[Cat.scala 29:58]
  wire [7:0] _GEN_88 = 8'h58 == _T_7[7:0] ? 8'h0 : _GEN_87; // @[Cat.scala 29:58]
  wire [7:0] _GEN_89 = 8'h59 == _T_7[7:0] ? 8'h0 : _GEN_88; // @[Cat.scala 29:58]
  wire [7:0] _GEN_90 = 8'h5a == _T_7[7:0] ? 8'h0 : _GEN_89; // @[Cat.scala 29:58]
  wire [7:0] _GEN_91 = 8'h5b == _T_7[7:0] ? 8'h0 : _GEN_90; // @[Cat.scala 29:58]
  wire [7:0] _GEN_92 = 8'h5c == _T_7[7:0] ? 8'h0 : _GEN_91; // @[Cat.scala 29:58]
  wire [7:0] _GEN_93 = 8'h5d == _T_7[7:0] ? 8'h0 : _GEN_92; // @[Cat.scala 29:58]
  wire [7:0] _GEN_94 = 8'h5e == _T_7[7:0] ? 8'h0 : _GEN_93; // @[Cat.scala 29:58]
  wire [7:0] _GEN_95 = 8'h5f == _T_7[7:0] ? 8'h0 : _GEN_94; // @[Cat.scala 29:58]
  wire [7:0] _GEN_96 = 8'h60 == _T_7[7:0] ? 8'h0 : _GEN_95; // @[Cat.scala 29:58]
  wire [7:0] _GEN_97 = 8'h61 == _T_7[7:0] ? 8'h0 : _GEN_96; // @[Cat.scala 29:58]
  wire [7:0] _GEN_98 = 8'h62 == _T_7[7:0] ? 8'h0 : _GEN_97; // @[Cat.scala 29:58]
  wire [7:0] _GEN_99 = 8'h63 == _T_7[7:0] ? 8'h0 : _GEN_98; // @[Cat.scala 29:58]
  wire [7:0] _GEN_100 = 8'h64 == _T_7[7:0] ? 8'h0 : _GEN_99; // @[Cat.scala 29:58]
  wire [7:0] _GEN_101 = 8'h65 == _T_7[7:0] ? 8'h0 : _GEN_100; // @[Cat.scala 29:58]
  wire [7:0] _GEN_102 = 8'h66 == _T_7[7:0] ? 8'h0 : _GEN_101; // @[Cat.scala 29:58]
  wire [7:0] _GEN_103 = 8'h67 == _T_7[7:0] ? 8'h0 : _GEN_102; // @[Cat.scala 29:58]
  wire [7:0] _GEN_104 = 8'h68 == _T_7[7:0] ? 8'h0 : _GEN_103; // @[Cat.scala 29:58]
  wire [7:0] _GEN_105 = 8'h69 == _T_7[7:0] ? 8'h0 : _GEN_104; // @[Cat.scala 29:58]
  wire [7:0] _GEN_106 = 8'h6a == _T_7[7:0] ? 8'h0 : _GEN_105; // @[Cat.scala 29:58]
  wire [7:0] _GEN_107 = 8'h6b == _T_7[7:0] ? 8'h0 : _GEN_106; // @[Cat.scala 29:58]
  wire [7:0] _GEN_108 = 8'h6c == _T_7[7:0] ? 8'h0 : _GEN_107; // @[Cat.scala 29:58]
  wire [7:0] _GEN_109 = 8'h6d == _T_7[7:0] ? 8'h0 : _GEN_108; // @[Cat.scala 29:58]
  wire [7:0] _GEN_110 = 8'h6e == _T_7[7:0] ? 8'h0 : _GEN_109; // @[Cat.scala 29:58]
  wire [7:0] _GEN_111 = 8'h6f == _T_7[7:0] ? 8'h0 : _GEN_110; // @[Cat.scala 29:58]
  wire [7:0] _GEN_112 = 8'h70 == _T_7[7:0] ? 8'h0 : _GEN_111; // @[Cat.scala 29:58]
  wire [7:0] _GEN_113 = 8'h71 == _T_7[7:0] ? 8'h0 : _GEN_112; // @[Cat.scala 29:58]
  wire [7:0] _GEN_114 = 8'h72 == _T_7[7:0] ? 8'h0 : _GEN_113; // @[Cat.scala 29:58]
  wire [7:0] _GEN_115 = 8'h73 == _T_7[7:0] ? 8'h0 : _GEN_114; // @[Cat.scala 29:58]
  wire [7:0] _GEN_116 = 8'h74 == _T_7[7:0] ? 8'h0 : _GEN_115; // @[Cat.scala 29:58]
  wire [7:0] _GEN_117 = 8'h75 == _T_7[7:0] ? 8'h0 : _GEN_116; // @[Cat.scala 29:58]
  wire [7:0] _GEN_118 = 8'h76 == _T_7[7:0] ? 8'h0 : _GEN_117; // @[Cat.scala 29:58]
  wire [7:0] _GEN_119 = 8'h77 == _T_7[7:0] ? 8'h0 : _GEN_118; // @[Cat.scala 29:58]
  wire [7:0] _GEN_120 = 8'h78 == _T_7[7:0] ? 8'h0 : _GEN_119; // @[Cat.scala 29:58]
  wire [7:0] _GEN_121 = 8'h79 == _T_7[7:0] ? 8'h0 : _GEN_120; // @[Cat.scala 29:58]
  wire [7:0] _GEN_122 = 8'h7a == _T_7[7:0] ? 8'h0 : _GEN_121; // @[Cat.scala 29:58]
  wire [7:0] _GEN_123 = 8'h7b == _T_7[7:0] ? 8'h0 : _GEN_122; // @[Cat.scala 29:58]
  wire [7:0] _GEN_124 = 8'h7c == _T_7[7:0] ? 8'h0 : _GEN_123; // @[Cat.scala 29:58]
  wire [7:0] _GEN_125 = 8'h7d == _T_7[7:0] ? 8'h0 : _GEN_124; // @[Cat.scala 29:58]
  wire [7:0] _GEN_126 = 8'h7e == _T_7[7:0] ? 8'h0 : _GEN_125; // @[Cat.scala 29:58]
  wire [7:0] _GEN_127 = 8'h7f == _T_7[7:0] ? 8'h0 : _GEN_126; // @[Cat.scala 29:58]
  wire [7:0] _GEN_128 = 8'h80 == _T_7[7:0] ? 8'h0 : _GEN_127; // @[Cat.scala 29:58]
  wire [7:0] _GEN_129 = 8'h81 == _T_7[7:0] ? 8'h0 : _GEN_128; // @[Cat.scala 29:58]
  wire [7:0] _GEN_130 = 8'h82 == _T_7[7:0] ? 8'h0 : _GEN_129; // @[Cat.scala 29:58]
  wire [7:0] _GEN_131 = 8'h83 == _T_7[7:0] ? 8'h0 : _GEN_130; // @[Cat.scala 29:58]
  wire [7:0] _GEN_132 = 8'h84 == _T_7[7:0] ? 8'h0 : _GEN_131; // @[Cat.scala 29:58]
  wire [7:0] _GEN_133 = 8'h85 == _T_7[7:0] ? 8'h0 : _GEN_132; // @[Cat.scala 29:58]
  wire [7:0] _GEN_134 = 8'h86 == _T_7[7:0] ? 8'h0 : _GEN_133; // @[Cat.scala 29:58]
  wire [7:0] _GEN_135 = 8'h87 == _T_7[7:0] ? 8'h0 : _GEN_134; // @[Cat.scala 29:58]
  wire [7:0] _GEN_136 = 8'h88 == _T_7[7:0] ? 8'h0 : _GEN_135; // @[Cat.scala 29:58]
  wire [7:0] _GEN_137 = 8'h89 == _T_7[7:0] ? 8'h0 : _GEN_136; // @[Cat.scala 29:58]
  wire [7:0] _GEN_138 = 8'h8a == _T_7[7:0] ? 8'h0 : _GEN_137; // @[Cat.scala 29:58]
  wire [7:0] _GEN_139 = 8'h8b == _T_7[7:0] ? 8'h0 : _GEN_138; // @[Cat.scala 29:58]
  wire [7:0] _GEN_140 = 8'h8c == _T_7[7:0] ? 8'h0 : _GEN_139; // @[Cat.scala 29:58]
  wire [7:0] _GEN_141 = 8'h8d == _T_7[7:0] ? 8'h0 : _GEN_140; // @[Cat.scala 29:58]
  wire [7:0] _GEN_142 = 8'h8e == _T_7[7:0] ? 8'h0 : _GEN_141; // @[Cat.scala 29:58]
  wire [7:0] _GEN_143 = 8'h8f == _T_7[7:0] ? 8'h0 : _GEN_142; // @[Cat.scala 29:58]
  wire [7:0] _GEN_144 = 8'h90 == _T_7[7:0] ? 8'h0 : _GEN_143; // @[Cat.scala 29:58]
  wire [7:0] _GEN_145 = 8'h91 == _T_7[7:0] ? 8'h0 : _GEN_144; // @[Cat.scala 29:58]
  wire [7:0] _GEN_146 = 8'h92 == _T_7[7:0] ? 8'h0 : _GEN_145; // @[Cat.scala 29:58]
  wire [7:0] _GEN_147 = 8'h93 == _T_7[7:0] ? 8'h0 : _GEN_146; // @[Cat.scala 29:58]
  wire [7:0] _GEN_148 = 8'h94 == _T_7[7:0] ? 8'h0 : _GEN_147; // @[Cat.scala 29:58]
  wire [7:0] _GEN_149 = 8'h95 == _T_7[7:0] ? 8'h0 : _GEN_148; // @[Cat.scala 29:58]
  wire [7:0] _GEN_150 = 8'h96 == _T_7[7:0] ? 8'h0 : _GEN_149; // @[Cat.scala 29:58]
  wire [7:0] _GEN_151 = 8'h97 == _T_7[7:0] ? 8'h0 : _GEN_150; // @[Cat.scala 29:58]
  wire [7:0] _GEN_152 = 8'h98 == _T_7[7:0] ? 8'h0 : _GEN_151; // @[Cat.scala 29:58]
  wire [7:0] _GEN_153 = 8'h99 == _T_7[7:0] ? 8'h0 : _GEN_152; // @[Cat.scala 29:58]
  wire [7:0] _GEN_154 = 8'h9a == _T_7[7:0] ? 8'h0 : _GEN_153; // @[Cat.scala 29:58]
  wire [7:0] _GEN_155 = 8'h9b == _T_7[7:0] ? 8'h0 : _GEN_154; // @[Cat.scala 29:58]
  wire [7:0] _GEN_156 = 8'h9c == _T_7[7:0] ? 8'h0 : _GEN_155; // @[Cat.scala 29:58]
  wire [7:0] _GEN_157 = 8'h9d == _T_7[7:0] ? 8'h0 : _GEN_156; // @[Cat.scala 29:58]
  wire [7:0] _GEN_158 = 8'h9e == _T_7[7:0] ? 8'h0 : _GEN_157; // @[Cat.scala 29:58]
  wire [7:0] _GEN_159 = 8'h9f == _T_7[7:0] ? 8'h0 : _GEN_158; // @[Cat.scala 29:58]
  wire [7:0] _GEN_160 = 8'ha0 == _T_7[7:0] ? 8'h0 : _GEN_159; // @[Cat.scala 29:58]
  wire [7:0] _GEN_161 = 8'ha1 == _T_7[7:0] ? 8'h0 : _GEN_160; // @[Cat.scala 29:58]
  wire [7:0] _GEN_162 = 8'ha2 == _T_7[7:0] ? 8'h0 : _GEN_161; // @[Cat.scala 29:58]
  wire [7:0] _GEN_163 = 8'ha3 == _T_7[7:0] ? 8'h0 : _GEN_162; // @[Cat.scala 29:58]
  wire [7:0] _GEN_164 = 8'ha4 == _T_7[7:0] ? 8'h0 : _GEN_163; // @[Cat.scala 29:58]
  wire [7:0] _GEN_165 = 8'ha5 == _T_7[7:0] ? 8'h0 : _GEN_164; // @[Cat.scala 29:58]
  wire [7:0] _GEN_166 = 8'ha6 == _T_7[7:0] ? 8'h0 : _GEN_165; // @[Cat.scala 29:58]
  wire [7:0] _GEN_167 = 8'ha7 == _T_7[7:0] ? 8'h0 : _GEN_166; // @[Cat.scala 29:58]
  wire [7:0] _GEN_168 = 8'ha8 == _T_7[7:0] ? 8'h0 : _GEN_167; // @[Cat.scala 29:58]
  wire [7:0] _GEN_169 = 8'ha9 == _T_7[7:0] ? 8'h0 : _GEN_168; // @[Cat.scala 29:58]
  wire [7:0] _GEN_170 = 8'haa == _T_7[7:0] ? 8'h0 : _GEN_169; // @[Cat.scala 29:58]
  wire [7:0] _GEN_171 = 8'hab == _T_7[7:0] ? 8'h0 : _GEN_170; // @[Cat.scala 29:58]
  wire [7:0] _GEN_172 = 8'hac == _T_7[7:0] ? 8'h0 : _GEN_171; // @[Cat.scala 29:58]
  wire [7:0] _GEN_173 = 8'had == _T_7[7:0] ? 8'h0 : _GEN_172; // @[Cat.scala 29:58]
  wire [7:0] _GEN_174 = 8'hae == _T_7[7:0] ? 8'h0 : _GEN_173; // @[Cat.scala 29:58]
  wire [7:0] _GEN_175 = 8'haf == _T_7[7:0] ? 8'h0 : _GEN_174; // @[Cat.scala 29:58]
  wire [7:0] _GEN_176 = 8'hb0 == _T_7[7:0] ? 8'h0 : _GEN_175; // @[Cat.scala 29:58]
  wire [7:0] _GEN_177 = 8'hb1 == _T_7[7:0] ? 8'h0 : _GEN_176; // @[Cat.scala 29:58]
  wire [7:0] _GEN_178 = 8'hb2 == _T_7[7:0] ? 8'h0 : _GEN_177; // @[Cat.scala 29:58]
  wire [7:0] _GEN_179 = 8'hb3 == _T_7[7:0] ? 8'h0 : _GEN_178; // @[Cat.scala 29:58]
  wire [7:0] _GEN_180 = 8'hb4 == _T_7[7:0] ? 8'h0 : _GEN_179; // @[Cat.scala 29:58]
  wire [7:0] _GEN_181 = 8'hb5 == _T_7[7:0] ? 8'h0 : _GEN_180; // @[Cat.scala 29:58]
  wire [7:0] _GEN_182 = 8'hb6 == _T_7[7:0] ? 8'h0 : _GEN_181; // @[Cat.scala 29:58]
  wire [7:0] _GEN_183 = 8'hb7 == _T_7[7:0] ? 8'h0 : _GEN_182; // @[Cat.scala 29:58]
  wire [7:0] _GEN_184 = 8'hb8 == _T_7[7:0] ? 8'h0 : _GEN_183; // @[Cat.scala 29:58]
  wire [7:0] _GEN_185 = 8'hb9 == _T_7[7:0] ? 8'h0 : _GEN_184; // @[Cat.scala 29:58]
  wire [7:0] _GEN_186 = 8'hba == _T_7[7:0] ? 8'h0 : _GEN_185; // @[Cat.scala 29:58]
  wire [7:0] _GEN_187 = 8'hbb == _T_7[7:0] ? 8'h0 : _GEN_186; // @[Cat.scala 29:58]
  wire [7:0] _GEN_188 = 8'hbc == _T_7[7:0] ? 8'h0 : _GEN_187; // @[Cat.scala 29:58]
  wire [7:0] _GEN_189 = 8'hbd == _T_7[7:0] ? 8'h0 : _GEN_188; // @[Cat.scala 29:58]
  wire [7:0] _GEN_190 = 8'hbe == _T_7[7:0] ? 8'h0 : _GEN_189; // @[Cat.scala 29:58]
  wire [7:0] _GEN_191 = 8'hbf == _T_7[7:0] ? 8'h0 : _GEN_190; // @[Cat.scala 29:58]
  wire [7:0] _GEN_192 = 8'hc0 == _T_7[7:0] ? 8'h0 : _GEN_191; // @[Cat.scala 29:58]
  wire [7:0] _GEN_193 = 8'hc1 == _T_7[7:0] ? 8'h0 : _GEN_192; // @[Cat.scala 29:58]
  wire [7:0] _GEN_194 = 8'hc2 == _T_7[7:0] ? 8'h0 : _GEN_193; // @[Cat.scala 29:58]
  wire [7:0] _GEN_195 = 8'hc3 == _T_7[7:0] ? 8'h0 : _GEN_194; // @[Cat.scala 29:58]
  wire [7:0] _GEN_196 = 8'hc4 == _T_7[7:0] ? 8'h0 : _GEN_195; // @[Cat.scala 29:58]
  wire [7:0] _GEN_197 = 8'hc5 == _T_7[7:0] ? 8'h0 : _GEN_196; // @[Cat.scala 29:58]
  wire [7:0] _GEN_198 = 8'hc6 == _T_7[7:0] ? 8'h0 : _GEN_197; // @[Cat.scala 29:58]
  wire [7:0] _GEN_199 = 8'hc7 == _T_7[7:0] ? 8'h0 : _GEN_198; // @[Cat.scala 29:58]
  wire [7:0] _GEN_200 = 8'hc8 == _T_7[7:0] ? 8'h0 : _GEN_199; // @[Cat.scala 29:58]
  wire [7:0] _GEN_201 = 8'hc9 == _T_7[7:0] ? 8'h0 : _GEN_200; // @[Cat.scala 29:58]
  wire [7:0] _GEN_202 = 8'hca == _T_7[7:0] ? 8'h0 : _GEN_201; // @[Cat.scala 29:58]
  wire [7:0] _GEN_203 = 8'hcb == _T_7[7:0] ? 8'h0 : _GEN_202; // @[Cat.scala 29:58]
  wire [7:0] _GEN_204 = 8'hcc == _T_7[7:0] ? 8'h0 : _GEN_203; // @[Cat.scala 29:58]
  wire [7:0] _GEN_205 = 8'hcd == _T_7[7:0] ? 8'h0 : _GEN_204; // @[Cat.scala 29:58]
  wire [7:0] _GEN_206 = 8'hce == _T_7[7:0] ? 8'h0 : _GEN_205; // @[Cat.scala 29:58]
  wire [7:0] _GEN_207 = 8'hcf == _T_7[7:0] ? 8'h0 : _GEN_206; // @[Cat.scala 29:58]
  wire [7:0] _GEN_208 = 8'hd0 == _T_7[7:0] ? 8'h0 : _GEN_207; // @[Cat.scala 29:58]
  wire [7:0] _GEN_209 = 8'hd1 == _T_7[7:0] ? 8'h0 : _GEN_208; // @[Cat.scala 29:58]
  wire [7:0] _GEN_210 = 8'hd2 == _T_7[7:0] ? 8'h0 : _GEN_209; // @[Cat.scala 29:58]
  wire [7:0] _GEN_211 = 8'hd3 == _T_7[7:0] ? 8'h0 : _GEN_210; // @[Cat.scala 29:58]
  wire [7:0] _GEN_212 = 8'hd4 == _T_7[7:0] ? 8'h0 : _GEN_211; // @[Cat.scala 29:58]
  wire [7:0] _GEN_213 = 8'hd5 == _T_7[7:0] ? 8'h0 : _GEN_212; // @[Cat.scala 29:58]
  wire [7:0] _GEN_214 = 8'hd6 == _T_7[7:0] ? 8'h0 : _GEN_213; // @[Cat.scala 29:58]
  wire [7:0] _GEN_215 = 8'hd7 == _T_7[7:0] ? 8'h0 : _GEN_214; // @[Cat.scala 29:58]
  wire [7:0] _GEN_216 = 8'hd8 == _T_7[7:0] ? 8'h0 : _GEN_215; // @[Cat.scala 29:58]
  wire [7:0] _GEN_217 = 8'hd9 == _T_7[7:0] ? 8'h0 : _GEN_216; // @[Cat.scala 29:58]
  wire [7:0] _GEN_218 = 8'hda == _T_7[7:0] ? 8'h0 : _GEN_217; // @[Cat.scala 29:58]
  wire [7:0] _GEN_219 = 8'hdb == _T_7[7:0] ? 8'h0 : _GEN_218; // @[Cat.scala 29:58]
  wire [7:0] _GEN_221 = 8'h1 == instrBus_pc[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_222 = 8'h2 == instrBus_pc[7:0] ? 8'h0 : _GEN_221; // @[Cat.scala 29:58]
  wire [7:0] _GEN_223 = 8'h3 == instrBus_pc[7:0] ? 8'hfe : _GEN_222; // @[Cat.scala 29:58]
  wire [7:0] _GEN_224 = 8'h4 == instrBus_pc[7:0] ? 8'h93 : _GEN_223; // @[Cat.scala 29:58]
  wire [7:0] _GEN_225 = 8'h5 == instrBus_pc[7:0] ? 8'h5 : _GEN_224; // @[Cat.scala 29:58]
  wire [7:0] _GEN_226 = 8'h6 == instrBus_pc[7:0] ? 8'h0 : _GEN_225; // @[Cat.scala 29:58]
  wire [7:0] _GEN_227 = 8'h7 == instrBus_pc[7:0] ? 8'hfc : _GEN_226; // @[Cat.scala 29:58]
  wire [7:0] _GEN_228 = 8'h8 == instrBus_pc[7:0] ? 8'h33 : _GEN_227; // @[Cat.scala 29:58]
  wire [7:0] _GEN_229 = 8'h9 == instrBus_pc[7:0] ? 8'h6 : _GEN_228; // @[Cat.scala 29:58]
  wire [7:0] _GEN_230 = 8'ha == instrBus_pc[7:0] ? 8'hb5 : _GEN_229; // @[Cat.scala 29:58]
  wire [7:0] _GEN_231 = 8'hb == instrBus_pc[7:0] ? 8'h0 : _GEN_230; // @[Cat.scala 29:58]
  wire [7:0] _GEN_232 = 8'hc == instrBus_pc[7:0] ? 8'h13 : _GEN_231; // @[Cat.scala 29:58]
  wire [7:0] _GEN_233 = 8'hd == instrBus_pc[7:0] ? 8'h5 : _GEN_232; // @[Cat.scala 29:58]
  wire [7:0] _GEN_234 = 8'he == instrBus_pc[7:0] ? 8'ha0 : _GEN_233; // @[Cat.scala 29:58]
  wire [7:0] _GEN_235 = 8'hf == instrBus_pc[7:0] ? 8'h0 : _GEN_234; // @[Cat.scala 29:58]
  wire [7:0] _GEN_236 = 8'h10 == instrBus_pc[7:0] ? 8'h73 : _GEN_235; // @[Cat.scala 29:58]
  wire [7:0] _GEN_237 = 8'h11 == instrBus_pc[7:0] ? 8'h0 : _GEN_236; // @[Cat.scala 29:58]
  wire [7:0] _GEN_238 = 8'h12 == instrBus_pc[7:0] ? 8'h0 : _GEN_237; // @[Cat.scala 29:58]
  wire [7:0] _GEN_239 = 8'h13 == instrBus_pc[7:0] ? 8'h0 : _GEN_238; // @[Cat.scala 29:58]
  wire [7:0] _GEN_240 = 8'h14 == instrBus_pc[7:0] ? 8'h0 : _GEN_239; // @[Cat.scala 29:58]
  wire [7:0] _GEN_241 = 8'h15 == instrBus_pc[7:0] ? 8'h0 : _GEN_240; // @[Cat.scala 29:58]
  wire [7:0] _GEN_242 = 8'h16 == instrBus_pc[7:0] ? 8'h0 : _GEN_241; // @[Cat.scala 29:58]
  wire [7:0] _GEN_243 = 8'h17 == instrBus_pc[7:0] ? 8'h0 : _GEN_242; // @[Cat.scala 29:58]
  wire [7:0] _GEN_244 = 8'h18 == instrBus_pc[7:0] ? 8'h0 : _GEN_243; // @[Cat.scala 29:58]
  wire [7:0] _GEN_245 = 8'h19 == instrBus_pc[7:0] ? 8'h0 : _GEN_244; // @[Cat.scala 29:58]
  wire [7:0] _GEN_246 = 8'h1a == instrBus_pc[7:0] ? 8'h0 : _GEN_245; // @[Cat.scala 29:58]
  wire [7:0] _GEN_247 = 8'h1b == instrBus_pc[7:0] ? 8'h0 : _GEN_246; // @[Cat.scala 29:58]
  wire [7:0] _GEN_248 = 8'h1c == instrBus_pc[7:0] ? 8'h0 : _GEN_247; // @[Cat.scala 29:58]
  wire [7:0] _GEN_249 = 8'h1d == instrBus_pc[7:0] ? 8'h0 : _GEN_248; // @[Cat.scala 29:58]
  wire [7:0] _GEN_250 = 8'h1e == instrBus_pc[7:0] ? 8'h0 : _GEN_249; // @[Cat.scala 29:58]
  wire [7:0] _GEN_251 = 8'h1f == instrBus_pc[7:0] ? 8'h0 : _GEN_250; // @[Cat.scala 29:58]
  wire [7:0] _GEN_252 = 8'h20 == instrBus_pc[7:0] ? 8'h0 : _GEN_251; // @[Cat.scala 29:58]
  wire [7:0] _GEN_253 = 8'h21 == instrBus_pc[7:0] ? 8'h0 : _GEN_252; // @[Cat.scala 29:58]
  wire [7:0] _GEN_254 = 8'h22 == instrBus_pc[7:0] ? 8'h0 : _GEN_253; // @[Cat.scala 29:58]
  wire [7:0] _GEN_255 = 8'h23 == instrBus_pc[7:0] ? 8'h0 : _GEN_254; // @[Cat.scala 29:58]
  wire [7:0] _GEN_256 = 8'h24 == instrBus_pc[7:0] ? 8'h0 : _GEN_255; // @[Cat.scala 29:58]
  wire [7:0] _GEN_257 = 8'h25 == instrBus_pc[7:0] ? 8'h0 : _GEN_256; // @[Cat.scala 29:58]
  wire [7:0] _GEN_258 = 8'h26 == instrBus_pc[7:0] ? 8'h0 : _GEN_257; // @[Cat.scala 29:58]
  wire [7:0] _GEN_259 = 8'h27 == instrBus_pc[7:0] ? 8'h0 : _GEN_258; // @[Cat.scala 29:58]
  wire [7:0] _GEN_260 = 8'h28 == instrBus_pc[7:0] ? 8'h0 : _GEN_259; // @[Cat.scala 29:58]
  wire [7:0] _GEN_261 = 8'h29 == instrBus_pc[7:0] ? 8'h0 : _GEN_260; // @[Cat.scala 29:58]
  wire [7:0] _GEN_262 = 8'h2a == instrBus_pc[7:0] ? 8'h0 : _GEN_261; // @[Cat.scala 29:58]
  wire [7:0] _GEN_263 = 8'h2b == instrBus_pc[7:0] ? 8'h0 : _GEN_262; // @[Cat.scala 29:58]
  wire [7:0] _GEN_264 = 8'h2c == instrBus_pc[7:0] ? 8'h0 : _GEN_263; // @[Cat.scala 29:58]
  wire [7:0] _GEN_265 = 8'h2d == instrBus_pc[7:0] ? 8'h0 : _GEN_264; // @[Cat.scala 29:58]
  wire [7:0] _GEN_266 = 8'h2e == instrBus_pc[7:0] ? 8'h0 : _GEN_265; // @[Cat.scala 29:58]
  wire [7:0] _GEN_267 = 8'h2f == instrBus_pc[7:0] ? 8'h0 : _GEN_266; // @[Cat.scala 29:58]
  wire [7:0] _GEN_268 = 8'h30 == instrBus_pc[7:0] ? 8'h0 : _GEN_267; // @[Cat.scala 29:58]
  wire [7:0] _GEN_269 = 8'h31 == instrBus_pc[7:0] ? 8'h0 : _GEN_268; // @[Cat.scala 29:58]
  wire [7:0] _GEN_270 = 8'h32 == instrBus_pc[7:0] ? 8'h0 : _GEN_269; // @[Cat.scala 29:58]
  wire [7:0] _GEN_271 = 8'h33 == instrBus_pc[7:0] ? 8'h0 : _GEN_270; // @[Cat.scala 29:58]
  wire [7:0] _GEN_272 = 8'h34 == instrBus_pc[7:0] ? 8'h0 : _GEN_271; // @[Cat.scala 29:58]
  wire [7:0] _GEN_273 = 8'h35 == instrBus_pc[7:0] ? 8'h0 : _GEN_272; // @[Cat.scala 29:58]
  wire [7:0] _GEN_274 = 8'h36 == instrBus_pc[7:0] ? 8'h0 : _GEN_273; // @[Cat.scala 29:58]
  wire [7:0] _GEN_275 = 8'h37 == instrBus_pc[7:0] ? 8'h0 : _GEN_274; // @[Cat.scala 29:58]
  wire [7:0] _GEN_276 = 8'h38 == instrBus_pc[7:0] ? 8'h0 : _GEN_275; // @[Cat.scala 29:58]
  wire [7:0] _GEN_277 = 8'h39 == instrBus_pc[7:0] ? 8'h0 : _GEN_276; // @[Cat.scala 29:58]
  wire [7:0] _GEN_278 = 8'h3a == instrBus_pc[7:0] ? 8'h0 : _GEN_277; // @[Cat.scala 29:58]
  wire [7:0] _GEN_279 = 8'h3b == instrBus_pc[7:0] ? 8'h0 : _GEN_278; // @[Cat.scala 29:58]
  wire [7:0] _GEN_280 = 8'h3c == instrBus_pc[7:0] ? 8'h0 : _GEN_279; // @[Cat.scala 29:58]
  wire [7:0] _GEN_281 = 8'h3d == instrBus_pc[7:0] ? 8'h0 : _GEN_280; // @[Cat.scala 29:58]
  wire [7:0] _GEN_282 = 8'h3e == instrBus_pc[7:0] ? 8'h0 : _GEN_281; // @[Cat.scala 29:58]
  wire [7:0] _GEN_283 = 8'h3f == instrBus_pc[7:0] ? 8'h0 : _GEN_282; // @[Cat.scala 29:58]
  wire [7:0] _GEN_284 = 8'h40 == instrBus_pc[7:0] ? 8'h0 : _GEN_283; // @[Cat.scala 29:58]
  wire [7:0] _GEN_285 = 8'h41 == instrBus_pc[7:0] ? 8'h0 : _GEN_284; // @[Cat.scala 29:58]
  wire [7:0] _GEN_286 = 8'h42 == instrBus_pc[7:0] ? 8'h0 : _GEN_285; // @[Cat.scala 29:58]
  wire [7:0] _GEN_287 = 8'h43 == instrBus_pc[7:0] ? 8'h0 : _GEN_286; // @[Cat.scala 29:58]
  wire [7:0] _GEN_288 = 8'h44 == instrBus_pc[7:0] ? 8'h0 : _GEN_287; // @[Cat.scala 29:58]
  wire [7:0] _GEN_289 = 8'h45 == instrBus_pc[7:0] ? 8'h0 : _GEN_288; // @[Cat.scala 29:58]
  wire [7:0] _GEN_290 = 8'h46 == instrBus_pc[7:0] ? 8'h0 : _GEN_289; // @[Cat.scala 29:58]
  wire [7:0] _GEN_291 = 8'h47 == instrBus_pc[7:0] ? 8'h0 : _GEN_290; // @[Cat.scala 29:58]
  wire [7:0] _GEN_292 = 8'h48 == instrBus_pc[7:0] ? 8'h0 : _GEN_291; // @[Cat.scala 29:58]
  wire [7:0] _GEN_293 = 8'h49 == instrBus_pc[7:0] ? 8'h0 : _GEN_292; // @[Cat.scala 29:58]
  wire [7:0] _GEN_294 = 8'h4a == instrBus_pc[7:0] ? 8'h0 : _GEN_293; // @[Cat.scala 29:58]
  wire [7:0] _GEN_295 = 8'h4b == instrBus_pc[7:0] ? 8'h0 : _GEN_294; // @[Cat.scala 29:58]
  wire [7:0] _GEN_296 = 8'h4c == instrBus_pc[7:0] ? 8'h0 : _GEN_295; // @[Cat.scala 29:58]
  wire [7:0] _GEN_297 = 8'h4d == instrBus_pc[7:0] ? 8'h0 : _GEN_296; // @[Cat.scala 29:58]
  wire [7:0] _GEN_298 = 8'h4e == instrBus_pc[7:0] ? 8'h0 : _GEN_297; // @[Cat.scala 29:58]
  wire [7:0] _GEN_299 = 8'h4f == instrBus_pc[7:0] ? 8'h0 : _GEN_298; // @[Cat.scala 29:58]
  wire [7:0] _GEN_300 = 8'h50 == instrBus_pc[7:0] ? 8'h0 : _GEN_299; // @[Cat.scala 29:58]
  wire [7:0] _GEN_301 = 8'h51 == instrBus_pc[7:0] ? 8'h0 : _GEN_300; // @[Cat.scala 29:58]
  wire [7:0] _GEN_302 = 8'h52 == instrBus_pc[7:0] ? 8'h0 : _GEN_301; // @[Cat.scala 29:58]
  wire [7:0] _GEN_303 = 8'h53 == instrBus_pc[7:0] ? 8'h0 : _GEN_302; // @[Cat.scala 29:58]
  wire [7:0] _GEN_304 = 8'h54 == instrBus_pc[7:0] ? 8'h0 : _GEN_303; // @[Cat.scala 29:58]
  wire [7:0] _GEN_305 = 8'h55 == instrBus_pc[7:0] ? 8'h0 : _GEN_304; // @[Cat.scala 29:58]
  wire [7:0] _GEN_306 = 8'h56 == instrBus_pc[7:0] ? 8'h0 : _GEN_305; // @[Cat.scala 29:58]
  wire [7:0] _GEN_307 = 8'h57 == instrBus_pc[7:0] ? 8'h0 : _GEN_306; // @[Cat.scala 29:58]
  wire [7:0] _GEN_308 = 8'h58 == instrBus_pc[7:0] ? 8'h0 : _GEN_307; // @[Cat.scala 29:58]
  wire [7:0] _GEN_309 = 8'h59 == instrBus_pc[7:0] ? 8'h0 : _GEN_308; // @[Cat.scala 29:58]
  wire [7:0] _GEN_310 = 8'h5a == instrBus_pc[7:0] ? 8'h0 : _GEN_309; // @[Cat.scala 29:58]
  wire [7:0] _GEN_311 = 8'h5b == instrBus_pc[7:0] ? 8'h0 : _GEN_310; // @[Cat.scala 29:58]
  wire [7:0] _GEN_312 = 8'h5c == instrBus_pc[7:0] ? 8'h0 : _GEN_311; // @[Cat.scala 29:58]
  wire [7:0] _GEN_313 = 8'h5d == instrBus_pc[7:0] ? 8'h0 : _GEN_312; // @[Cat.scala 29:58]
  wire [7:0] _GEN_314 = 8'h5e == instrBus_pc[7:0] ? 8'h0 : _GEN_313; // @[Cat.scala 29:58]
  wire [7:0] _GEN_315 = 8'h5f == instrBus_pc[7:0] ? 8'h0 : _GEN_314; // @[Cat.scala 29:58]
  wire [7:0] _GEN_316 = 8'h60 == instrBus_pc[7:0] ? 8'h0 : _GEN_315; // @[Cat.scala 29:58]
  wire [7:0] _GEN_317 = 8'h61 == instrBus_pc[7:0] ? 8'h0 : _GEN_316; // @[Cat.scala 29:58]
  wire [7:0] _GEN_318 = 8'h62 == instrBus_pc[7:0] ? 8'h0 : _GEN_317; // @[Cat.scala 29:58]
  wire [7:0] _GEN_319 = 8'h63 == instrBus_pc[7:0] ? 8'h0 : _GEN_318; // @[Cat.scala 29:58]
  wire [7:0] _GEN_320 = 8'h64 == instrBus_pc[7:0] ? 8'h0 : _GEN_319; // @[Cat.scala 29:58]
  wire [7:0] _GEN_321 = 8'h65 == instrBus_pc[7:0] ? 8'h0 : _GEN_320; // @[Cat.scala 29:58]
  wire [7:0] _GEN_322 = 8'h66 == instrBus_pc[7:0] ? 8'h0 : _GEN_321; // @[Cat.scala 29:58]
  wire [7:0] _GEN_323 = 8'h67 == instrBus_pc[7:0] ? 8'h0 : _GEN_322; // @[Cat.scala 29:58]
  wire [7:0] _GEN_324 = 8'h68 == instrBus_pc[7:0] ? 8'h0 : _GEN_323; // @[Cat.scala 29:58]
  wire [7:0] _GEN_325 = 8'h69 == instrBus_pc[7:0] ? 8'h0 : _GEN_324; // @[Cat.scala 29:58]
  wire [7:0] _GEN_326 = 8'h6a == instrBus_pc[7:0] ? 8'h0 : _GEN_325; // @[Cat.scala 29:58]
  wire [7:0] _GEN_327 = 8'h6b == instrBus_pc[7:0] ? 8'h0 : _GEN_326; // @[Cat.scala 29:58]
  wire [7:0] _GEN_328 = 8'h6c == instrBus_pc[7:0] ? 8'h0 : _GEN_327; // @[Cat.scala 29:58]
  wire [7:0] _GEN_329 = 8'h6d == instrBus_pc[7:0] ? 8'h0 : _GEN_328; // @[Cat.scala 29:58]
  wire [7:0] _GEN_330 = 8'h6e == instrBus_pc[7:0] ? 8'h0 : _GEN_329; // @[Cat.scala 29:58]
  wire [7:0] _GEN_331 = 8'h6f == instrBus_pc[7:0] ? 8'h0 : _GEN_330; // @[Cat.scala 29:58]
  wire [7:0] _GEN_332 = 8'h70 == instrBus_pc[7:0] ? 8'h0 : _GEN_331; // @[Cat.scala 29:58]
  wire [7:0] _GEN_333 = 8'h71 == instrBus_pc[7:0] ? 8'h0 : _GEN_332; // @[Cat.scala 29:58]
  wire [7:0] _GEN_334 = 8'h72 == instrBus_pc[7:0] ? 8'h0 : _GEN_333; // @[Cat.scala 29:58]
  wire [7:0] _GEN_335 = 8'h73 == instrBus_pc[7:0] ? 8'h0 : _GEN_334; // @[Cat.scala 29:58]
  wire [7:0] _GEN_336 = 8'h74 == instrBus_pc[7:0] ? 8'h0 : _GEN_335; // @[Cat.scala 29:58]
  wire [7:0] _GEN_337 = 8'h75 == instrBus_pc[7:0] ? 8'h0 : _GEN_336; // @[Cat.scala 29:58]
  wire [7:0] _GEN_338 = 8'h76 == instrBus_pc[7:0] ? 8'h0 : _GEN_337; // @[Cat.scala 29:58]
  wire [7:0] _GEN_339 = 8'h77 == instrBus_pc[7:0] ? 8'h0 : _GEN_338; // @[Cat.scala 29:58]
  wire [7:0] _GEN_340 = 8'h78 == instrBus_pc[7:0] ? 8'h0 : _GEN_339; // @[Cat.scala 29:58]
  wire [7:0] _GEN_341 = 8'h79 == instrBus_pc[7:0] ? 8'h0 : _GEN_340; // @[Cat.scala 29:58]
  wire [7:0] _GEN_342 = 8'h7a == instrBus_pc[7:0] ? 8'h0 : _GEN_341; // @[Cat.scala 29:58]
  wire [7:0] _GEN_343 = 8'h7b == instrBus_pc[7:0] ? 8'h0 : _GEN_342; // @[Cat.scala 29:58]
  wire [7:0] _GEN_344 = 8'h7c == instrBus_pc[7:0] ? 8'h0 : _GEN_343; // @[Cat.scala 29:58]
  wire [7:0] _GEN_345 = 8'h7d == instrBus_pc[7:0] ? 8'h0 : _GEN_344; // @[Cat.scala 29:58]
  wire [7:0] _GEN_346 = 8'h7e == instrBus_pc[7:0] ? 8'h0 : _GEN_345; // @[Cat.scala 29:58]
  wire [7:0] _GEN_347 = 8'h7f == instrBus_pc[7:0] ? 8'h0 : _GEN_346; // @[Cat.scala 29:58]
  wire [7:0] _GEN_348 = 8'h80 == instrBus_pc[7:0] ? 8'h0 : _GEN_347; // @[Cat.scala 29:58]
  wire [7:0] _GEN_349 = 8'h81 == instrBus_pc[7:0] ? 8'h0 : _GEN_348; // @[Cat.scala 29:58]
  wire [7:0] _GEN_350 = 8'h82 == instrBus_pc[7:0] ? 8'h0 : _GEN_349; // @[Cat.scala 29:58]
  wire [7:0] _GEN_351 = 8'h83 == instrBus_pc[7:0] ? 8'h0 : _GEN_350; // @[Cat.scala 29:58]
  wire [7:0] _GEN_352 = 8'h84 == instrBus_pc[7:0] ? 8'h0 : _GEN_351; // @[Cat.scala 29:58]
  wire [7:0] _GEN_353 = 8'h85 == instrBus_pc[7:0] ? 8'h0 : _GEN_352; // @[Cat.scala 29:58]
  wire [7:0] _GEN_354 = 8'h86 == instrBus_pc[7:0] ? 8'h0 : _GEN_353; // @[Cat.scala 29:58]
  wire [7:0] _GEN_355 = 8'h87 == instrBus_pc[7:0] ? 8'h0 : _GEN_354; // @[Cat.scala 29:58]
  wire [7:0] _GEN_356 = 8'h88 == instrBus_pc[7:0] ? 8'h0 : _GEN_355; // @[Cat.scala 29:58]
  wire [7:0] _GEN_357 = 8'h89 == instrBus_pc[7:0] ? 8'h0 : _GEN_356; // @[Cat.scala 29:58]
  wire [7:0] _GEN_358 = 8'h8a == instrBus_pc[7:0] ? 8'h0 : _GEN_357; // @[Cat.scala 29:58]
  wire [7:0] _GEN_359 = 8'h8b == instrBus_pc[7:0] ? 8'h0 : _GEN_358; // @[Cat.scala 29:58]
  wire [7:0] _GEN_360 = 8'h8c == instrBus_pc[7:0] ? 8'h0 : _GEN_359; // @[Cat.scala 29:58]
  wire [7:0] _GEN_361 = 8'h8d == instrBus_pc[7:0] ? 8'h0 : _GEN_360; // @[Cat.scala 29:58]
  wire [7:0] _GEN_362 = 8'h8e == instrBus_pc[7:0] ? 8'h0 : _GEN_361; // @[Cat.scala 29:58]
  wire [7:0] _GEN_363 = 8'h8f == instrBus_pc[7:0] ? 8'h0 : _GEN_362; // @[Cat.scala 29:58]
  wire [7:0] _GEN_364 = 8'h90 == instrBus_pc[7:0] ? 8'h0 : _GEN_363; // @[Cat.scala 29:58]
  wire [7:0] _GEN_365 = 8'h91 == instrBus_pc[7:0] ? 8'h0 : _GEN_364; // @[Cat.scala 29:58]
  wire [7:0] _GEN_366 = 8'h92 == instrBus_pc[7:0] ? 8'h0 : _GEN_365; // @[Cat.scala 29:58]
  wire [7:0] _GEN_367 = 8'h93 == instrBus_pc[7:0] ? 8'h0 : _GEN_366; // @[Cat.scala 29:58]
  wire [7:0] _GEN_368 = 8'h94 == instrBus_pc[7:0] ? 8'h0 : _GEN_367; // @[Cat.scala 29:58]
  wire [7:0] _GEN_369 = 8'h95 == instrBus_pc[7:0] ? 8'h0 : _GEN_368; // @[Cat.scala 29:58]
  wire [7:0] _GEN_370 = 8'h96 == instrBus_pc[7:0] ? 8'h0 : _GEN_369; // @[Cat.scala 29:58]
  wire [7:0] _GEN_371 = 8'h97 == instrBus_pc[7:0] ? 8'h0 : _GEN_370; // @[Cat.scala 29:58]
  wire [7:0] _GEN_372 = 8'h98 == instrBus_pc[7:0] ? 8'h0 : _GEN_371; // @[Cat.scala 29:58]
  wire [7:0] _GEN_373 = 8'h99 == instrBus_pc[7:0] ? 8'h0 : _GEN_372; // @[Cat.scala 29:58]
  wire [7:0] _GEN_374 = 8'h9a == instrBus_pc[7:0] ? 8'h0 : _GEN_373; // @[Cat.scala 29:58]
  wire [7:0] _GEN_375 = 8'h9b == instrBus_pc[7:0] ? 8'h0 : _GEN_374; // @[Cat.scala 29:58]
  wire [7:0] _GEN_376 = 8'h9c == instrBus_pc[7:0] ? 8'h0 : _GEN_375; // @[Cat.scala 29:58]
  wire [7:0] _GEN_377 = 8'h9d == instrBus_pc[7:0] ? 8'h0 : _GEN_376; // @[Cat.scala 29:58]
  wire [7:0] _GEN_378 = 8'h9e == instrBus_pc[7:0] ? 8'h0 : _GEN_377; // @[Cat.scala 29:58]
  wire [7:0] _GEN_379 = 8'h9f == instrBus_pc[7:0] ? 8'h0 : _GEN_378; // @[Cat.scala 29:58]
  wire [7:0] _GEN_380 = 8'ha0 == instrBus_pc[7:0] ? 8'h0 : _GEN_379; // @[Cat.scala 29:58]
  wire [7:0] _GEN_381 = 8'ha1 == instrBus_pc[7:0] ? 8'h0 : _GEN_380; // @[Cat.scala 29:58]
  wire [7:0] _GEN_382 = 8'ha2 == instrBus_pc[7:0] ? 8'h0 : _GEN_381; // @[Cat.scala 29:58]
  wire [7:0] _GEN_383 = 8'ha3 == instrBus_pc[7:0] ? 8'h0 : _GEN_382; // @[Cat.scala 29:58]
  wire [7:0] _GEN_384 = 8'ha4 == instrBus_pc[7:0] ? 8'h0 : _GEN_383; // @[Cat.scala 29:58]
  wire [7:0] _GEN_385 = 8'ha5 == instrBus_pc[7:0] ? 8'h0 : _GEN_384; // @[Cat.scala 29:58]
  wire [7:0] _GEN_386 = 8'ha6 == instrBus_pc[7:0] ? 8'h0 : _GEN_385; // @[Cat.scala 29:58]
  wire [7:0] _GEN_387 = 8'ha7 == instrBus_pc[7:0] ? 8'h0 : _GEN_386; // @[Cat.scala 29:58]
  wire [7:0] _GEN_388 = 8'ha8 == instrBus_pc[7:0] ? 8'h0 : _GEN_387; // @[Cat.scala 29:58]
  wire [7:0] _GEN_389 = 8'ha9 == instrBus_pc[7:0] ? 8'h0 : _GEN_388; // @[Cat.scala 29:58]
  wire [7:0] _GEN_390 = 8'haa == instrBus_pc[7:0] ? 8'h0 : _GEN_389; // @[Cat.scala 29:58]
  wire [7:0] _GEN_391 = 8'hab == instrBus_pc[7:0] ? 8'h0 : _GEN_390; // @[Cat.scala 29:58]
  wire [7:0] _GEN_392 = 8'hac == instrBus_pc[7:0] ? 8'h0 : _GEN_391; // @[Cat.scala 29:58]
  wire [7:0] _GEN_393 = 8'had == instrBus_pc[7:0] ? 8'h0 : _GEN_392; // @[Cat.scala 29:58]
  wire [7:0] _GEN_394 = 8'hae == instrBus_pc[7:0] ? 8'h0 : _GEN_393; // @[Cat.scala 29:58]
  wire [7:0] _GEN_395 = 8'haf == instrBus_pc[7:0] ? 8'h0 : _GEN_394; // @[Cat.scala 29:58]
  wire [7:0] _GEN_396 = 8'hb0 == instrBus_pc[7:0] ? 8'h0 : _GEN_395; // @[Cat.scala 29:58]
  wire [7:0] _GEN_397 = 8'hb1 == instrBus_pc[7:0] ? 8'h0 : _GEN_396; // @[Cat.scala 29:58]
  wire [7:0] _GEN_398 = 8'hb2 == instrBus_pc[7:0] ? 8'h0 : _GEN_397; // @[Cat.scala 29:58]
  wire [7:0] _GEN_399 = 8'hb3 == instrBus_pc[7:0] ? 8'h0 : _GEN_398; // @[Cat.scala 29:58]
  wire [7:0] _GEN_400 = 8'hb4 == instrBus_pc[7:0] ? 8'h0 : _GEN_399; // @[Cat.scala 29:58]
  wire [7:0] _GEN_401 = 8'hb5 == instrBus_pc[7:0] ? 8'h0 : _GEN_400; // @[Cat.scala 29:58]
  wire [7:0] _GEN_402 = 8'hb6 == instrBus_pc[7:0] ? 8'h0 : _GEN_401; // @[Cat.scala 29:58]
  wire [7:0] _GEN_403 = 8'hb7 == instrBus_pc[7:0] ? 8'h0 : _GEN_402; // @[Cat.scala 29:58]
  wire [7:0] _GEN_404 = 8'hb8 == instrBus_pc[7:0] ? 8'h0 : _GEN_403; // @[Cat.scala 29:58]
  wire [7:0] _GEN_405 = 8'hb9 == instrBus_pc[7:0] ? 8'h0 : _GEN_404; // @[Cat.scala 29:58]
  wire [7:0] _GEN_406 = 8'hba == instrBus_pc[7:0] ? 8'h0 : _GEN_405; // @[Cat.scala 29:58]
  wire [7:0] _GEN_407 = 8'hbb == instrBus_pc[7:0] ? 8'h0 : _GEN_406; // @[Cat.scala 29:58]
  wire [7:0] _GEN_408 = 8'hbc == instrBus_pc[7:0] ? 8'h0 : _GEN_407; // @[Cat.scala 29:58]
  wire [7:0] _GEN_409 = 8'hbd == instrBus_pc[7:0] ? 8'h0 : _GEN_408; // @[Cat.scala 29:58]
  wire [7:0] _GEN_410 = 8'hbe == instrBus_pc[7:0] ? 8'h0 : _GEN_409; // @[Cat.scala 29:58]
  wire [7:0] _GEN_411 = 8'hbf == instrBus_pc[7:0] ? 8'h0 : _GEN_410; // @[Cat.scala 29:58]
  wire [7:0] _GEN_412 = 8'hc0 == instrBus_pc[7:0] ? 8'h0 : _GEN_411; // @[Cat.scala 29:58]
  wire [7:0] _GEN_413 = 8'hc1 == instrBus_pc[7:0] ? 8'h0 : _GEN_412; // @[Cat.scala 29:58]
  wire [7:0] _GEN_414 = 8'hc2 == instrBus_pc[7:0] ? 8'h0 : _GEN_413; // @[Cat.scala 29:58]
  wire [7:0] _GEN_415 = 8'hc3 == instrBus_pc[7:0] ? 8'h0 : _GEN_414; // @[Cat.scala 29:58]
  wire [7:0] _GEN_416 = 8'hc4 == instrBus_pc[7:0] ? 8'h0 : _GEN_415; // @[Cat.scala 29:58]
  wire [7:0] _GEN_417 = 8'hc5 == instrBus_pc[7:0] ? 8'h0 : _GEN_416; // @[Cat.scala 29:58]
  wire [7:0] _GEN_418 = 8'hc6 == instrBus_pc[7:0] ? 8'h0 : _GEN_417; // @[Cat.scala 29:58]
  wire [7:0] _GEN_419 = 8'hc7 == instrBus_pc[7:0] ? 8'h0 : _GEN_418; // @[Cat.scala 29:58]
  wire [7:0] _GEN_420 = 8'hc8 == instrBus_pc[7:0] ? 8'h0 : _GEN_419; // @[Cat.scala 29:58]
  wire [7:0] _GEN_421 = 8'hc9 == instrBus_pc[7:0] ? 8'h0 : _GEN_420; // @[Cat.scala 29:58]
  wire [7:0] _GEN_422 = 8'hca == instrBus_pc[7:0] ? 8'h0 : _GEN_421; // @[Cat.scala 29:58]
  wire [7:0] _GEN_423 = 8'hcb == instrBus_pc[7:0] ? 8'h0 : _GEN_422; // @[Cat.scala 29:58]
  wire [7:0] _GEN_424 = 8'hcc == instrBus_pc[7:0] ? 8'h0 : _GEN_423; // @[Cat.scala 29:58]
  wire [7:0] _GEN_425 = 8'hcd == instrBus_pc[7:0] ? 8'h0 : _GEN_424; // @[Cat.scala 29:58]
  wire [7:0] _GEN_426 = 8'hce == instrBus_pc[7:0] ? 8'h0 : _GEN_425; // @[Cat.scala 29:58]
  wire [7:0] _GEN_427 = 8'hcf == instrBus_pc[7:0] ? 8'h0 : _GEN_426; // @[Cat.scala 29:58]
  wire [7:0] _GEN_428 = 8'hd0 == instrBus_pc[7:0] ? 8'h0 : _GEN_427; // @[Cat.scala 29:58]
  wire [7:0] _GEN_429 = 8'hd1 == instrBus_pc[7:0] ? 8'h0 : _GEN_428; // @[Cat.scala 29:58]
  wire [7:0] _GEN_430 = 8'hd2 == instrBus_pc[7:0] ? 8'h0 : _GEN_429; // @[Cat.scala 29:58]
  wire [7:0] _GEN_431 = 8'hd3 == instrBus_pc[7:0] ? 8'h0 : _GEN_430; // @[Cat.scala 29:58]
  wire [7:0] _GEN_432 = 8'hd4 == instrBus_pc[7:0] ? 8'h0 : _GEN_431; // @[Cat.scala 29:58]
  wire [7:0] _GEN_433 = 8'hd5 == instrBus_pc[7:0] ? 8'h0 : _GEN_432; // @[Cat.scala 29:58]
  wire [7:0] _GEN_434 = 8'hd6 == instrBus_pc[7:0] ? 8'h0 : _GEN_433; // @[Cat.scala 29:58]
  wire [7:0] _GEN_435 = 8'hd7 == instrBus_pc[7:0] ? 8'h0 : _GEN_434; // @[Cat.scala 29:58]
  wire [7:0] _GEN_436 = 8'hd8 == instrBus_pc[7:0] ? 8'h0 : _GEN_435; // @[Cat.scala 29:58]
  wire [7:0] _GEN_437 = 8'hd9 == instrBus_pc[7:0] ? 8'h0 : _GEN_436; // @[Cat.scala 29:58]
  wire [7:0] _GEN_438 = 8'hda == instrBus_pc[7:0] ? 8'h0 : _GEN_437; // @[Cat.scala 29:58]
  wire [7:0] _GEN_439 = 8'hdb == instrBus_pc[7:0] ? 8'h0 : _GEN_438; // @[Cat.scala 29:58]
  wire [15:0] _T_10 = {_GEN_219,_GEN_439}; // @[Cat.scala 29:58]
  wire [7:0] _GEN_441 = 8'h1 == _T_1[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_442 = 8'h2 == _T_1[7:0] ? 8'h0 : _GEN_441; // @[Cat.scala 29:58]
  wire [7:0] _GEN_443 = 8'h3 == _T_1[7:0] ? 8'hfe : _GEN_442; // @[Cat.scala 29:58]
  wire [7:0] _GEN_444 = 8'h4 == _T_1[7:0] ? 8'h93 : _GEN_443; // @[Cat.scala 29:58]
  wire [7:0] _GEN_445 = 8'h5 == _T_1[7:0] ? 8'h5 : _GEN_444; // @[Cat.scala 29:58]
  wire [7:0] _GEN_446 = 8'h6 == _T_1[7:0] ? 8'h0 : _GEN_445; // @[Cat.scala 29:58]
  wire [7:0] _GEN_447 = 8'h7 == _T_1[7:0] ? 8'hfc : _GEN_446; // @[Cat.scala 29:58]
  wire [7:0] _GEN_448 = 8'h8 == _T_1[7:0] ? 8'h33 : _GEN_447; // @[Cat.scala 29:58]
  wire [7:0] _GEN_449 = 8'h9 == _T_1[7:0] ? 8'h6 : _GEN_448; // @[Cat.scala 29:58]
  wire [7:0] _GEN_450 = 8'ha == _T_1[7:0] ? 8'hb5 : _GEN_449; // @[Cat.scala 29:58]
  wire [7:0] _GEN_451 = 8'hb == _T_1[7:0] ? 8'h0 : _GEN_450; // @[Cat.scala 29:58]
  wire [7:0] _GEN_452 = 8'hc == _T_1[7:0] ? 8'h13 : _GEN_451; // @[Cat.scala 29:58]
  wire [7:0] _GEN_453 = 8'hd == _T_1[7:0] ? 8'h5 : _GEN_452; // @[Cat.scala 29:58]
  wire [7:0] _GEN_454 = 8'he == _T_1[7:0] ? 8'ha0 : _GEN_453; // @[Cat.scala 29:58]
  wire [7:0] _GEN_455 = 8'hf == _T_1[7:0] ? 8'h0 : _GEN_454; // @[Cat.scala 29:58]
  wire [7:0] _GEN_456 = 8'h10 == _T_1[7:0] ? 8'h73 : _GEN_455; // @[Cat.scala 29:58]
  wire [7:0] _GEN_457 = 8'h11 == _T_1[7:0] ? 8'h0 : _GEN_456; // @[Cat.scala 29:58]
  wire [7:0] _GEN_458 = 8'h12 == _T_1[7:0] ? 8'h0 : _GEN_457; // @[Cat.scala 29:58]
  wire [7:0] _GEN_459 = 8'h13 == _T_1[7:0] ? 8'h0 : _GEN_458; // @[Cat.scala 29:58]
  wire [7:0] _GEN_460 = 8'h14 == _T_1[7:0] ? 8'h0 : _GEN_459; // @[Cat.scala 29:58]
  wire [7:0] _GEN_461 = 8'h15 == _T_1[7:0] ? 8'h0 : _GEN_460; // @[Cat.scala 29:58]
  wire [7:0] _GEN_462 = 8'h16 == _T_1[7:0] ? 8'h0 : _GEN_461; // @[Cat.scala 29:58]
  wire [7:0] _GEN_463 = 8'h17 == _T_1[7:0] ? 8'h0 : _GEN_462; // @[Cat.scala 29:58]
  wire [7:0] _GEN_464 = 8'h18 == _T_1[7:0] ? 8'h0 : _GEN_463; // @[Cat.scala 29:58]
  wire [7:0] _GEN_465 = 8'h19 == _T_1[7:0] ? 8'h0 : _GEN_464; // @[Cat.scala 29:58]
  wire [7:0] _GEN_466 = 8'h1a == _T_1[7:0] ? 8'h0 : _GEN_465; // @[Cat.scala 29:58]
  wire [7:0] _GEN_467 = 8'h1b == _T_1[7:0] ? 8'h0 : _GEN_466; // @[Cat.scala 29:58]
  wire [7:0] _GEN_468 = 8'h1c == _T_1[7:0] ? 8'h0 : _GEN_467; // @[Cat.scala 29:58]
  wire [7:0] _GEN_469 = 8'h1d == _T_1[7:0] ? 8'h0 : _GEN_468; // @[Cat.scala 29:58]
  wire [7:0] _GEN_470 = 8'h1e == _T_1[7:0] ? 8'h0 : _GEN_469; // @[Cat.scala 29:58]
  wire [7:0] _GEN_471 = 8'h1f == _T_1[7:0] ? 8'h0 : _GEN_470; // @[Cat.scala 29:58]
  wire [7:0] _GEN_472 = 8'h20 == _T_1[7:0] ? 8'h0 : _GEN_471; // @[Cat.scala 29:58]
  wire [7:0] _GEN_473 = 8'h21 == _T_1[7:0] ? 8'h0 : _GEN_472; // @[Cat.scala 29:58]
  wire [7:0] _GEN_474 = 8'h22 == _T_1[7:0] ? 8'h0 : _GEN_473; // @[Cat.scala 29:58]
  wire [7:0] _GEN_475 = 8'h23 == _T_1[7:0] ? 8'h0 : _GEN_474; // @[Cat.scala 29:58]
  wire [7:0] _GEN_476 = 8'h24 == _T_1[7:0] ? 8'h0 : _GEN_475; // @[Cat.scala 29:58]
  wire [7:0] _GEN_477 = 8'h25 == _T_1[7:0] ? 8'h0 : _GEN_476; // @[Cat.scala 29:58]
  wire [7:0] _GEN_478 = 8'h26 == _T_1[7:0] ? 8'h0 : _GEN_477; // @[Cat.scala 29:58]
  wire [7:0] _GEN_479 = 8'h27 == _T_1[7:0] ? 8'h0 : _GEN_478; // @[Cat.scala 29:58]
  wire [7:0] _GEN_480 = 8'h28 == _T_1[7:0] ? 8'h0 : _GEN_479; // @[Cat.scala 29:58]
  wire [7:0] _GEN_481 = 8'h29 == _T_1[7:0] ? 8'h0 : _GEN_480; // @[Cat.scala 29:58]
  wire [7:0] _GEN_482 = 8'h2a == _T_1[7:0] ? 8'h0 : _GEN_481; // @[Cat.scala 29:58]
  wire [7:0] _GEN_483 = 8'h2b == _T_1[7:0] ? 8'h0 : _GEN_482; // @[Cat.scala 29:58]
  wire [7:0] _GEN_484 = 8'h2c == _T_1[7:0] ? 8'h0 : _GEN_483; // @[Cat.scala 29:58]
  wire [7:0] _GEN_485 = 8'h2d == _T_1[7:0] ? 8'h0 : _GEN_484; // @[Cat.scala 29:58]
  wire [7:0] _GEN_486 = 8'h2e == _T_1[7:0] ? 8'h0 : _GEN_485; // @[Cat.scala 29:58]
  wire [7:0] _GEN_487 = 8'h2f == _T_1[7:0] ? 8'h0 : _GEN_486; // @[Cat.scala 29:58]
  wire [7:0] _GEN_488 = 8'h30 == _T_1[7:0] ? 8'h0 : _GEN_487; // @[Cat.scala 29:58]
  wire [7:0] _GEN_489 = 8'h31 == _T_1[7:0] ? 8'h0 : _GEN_488; // @[Cat.scala 29:58]
  wire [7:0] _GEN_490 = 8'h32 == _T_1[7:0] ? 8'h0 : _GEN_489; // @[Cat.scala 29:58]
  wire [7:0] _GEN_491 = 8'h33 == _T_1[7:0] ? 8'h0 : _GEN_490; // @[Cat.scala 29:58]
  wire [7:0] _GEN_492 = 8'h34 == _T_1[7:0] ? 8'h0 : _GEN_491; // @[Cat.scala 29:58]
  wire [7:0] _GEN_493 = 8'h35 == _T_1[7:0] ? 8'h0 : _GEN_492; // @[Cat.scala 29:58]
  wire [7:0] _GEN_494 = 8'h36 == _T_1[7:0] ? 8'h0 : _GEN_493; // @[Cat.scala 29:58]
  wire [7:0] _GEN_495 = 8'h37 == _T_1[7:0] ? 8'h0 : _GEN_494; // @[Cat.scala 29:58]
  wire [7:0] _GEN_496 = 8'h38 == _T_1[7:0] ? 8'h0 : _GEN_495; // @[Cat.scala 29:58]
  wire [7:0] _GEN_497 = 8'h39 == _T_1[7:0] ? 8'h0 : _GEN_496; // @[Cat.scala 29:58]
  wire [7:0] _GEN_498 = 8'h3a == _T_1[7:0] ? 8'h0 : _GEN_497; // @[Cat.scala 29:58]
  wire [7:0] _GEN_499 = 8'h3b == _T_1[7:0] ? 8'h0 : _GEN_498; // @[Cat.scala 29:58]
  wire [7:0] _GEN_500 = 8'h3c == _T_1[7:0] ? 8'h0 : _GEN_499; // @[Cat.scala 29:58]
  wire [7:0] _GEN_501 = 8'h3d == _T_1[7:0] ? 8'h0 : _GEN_500; // @[Cat.scala 29:58]
  wire [7:0] _GEN_502 = 8'h3e == _T_1[7:0] ? 8'h0 : _GEN_501; // @[Cat.scala 29:58]
  wire [7:0] _GEN_503 = 8'h3f == _T_1[7:0] ? 8'h0 : _GEN_502; // @[Cat.scala 29:58]
  wire [7:0] _GEN_504 = 8'h40 == _T_1[7:0] ? 8'h0 : _GEN_503; // @[Cat.scala 29:58]
  wire [7:0] _GEN_505 = 8'h41 == _T_1[7:0] ? 8'h0 : _GEN_504; // @[Cat.scala 29:58]
  wire [7:0] _GEN_506 = 8'h42 == _T_1[7:0] ? 8'h0 : _GEN_505; // @[Cat.scala 29:58]
  wire [7:0] _GEN_507 = 8'h43 == _T_1[7:0] ? 8'h0 : _GEN_506; // @[Cat.scala 29:58]
  wire [7:0] _GEN_508 = 8'h44 == _T_1[7:0] ? 8'h0 : _GEN_507; // @[Cat.scala 29:58]
  wire [7:0] _GEN_509 = 8'h45 == _T_1[7:0] ? 8'h0 : _GEN_508; // @[Cat.scala 29:58]
  wire [7:0] _GEN_510 = 8'h46 == _T_1[7:0] ? 8'h0 : _GEN_509; // @[Cat.scala 29:58]
  wire [7:0] _GEN_511 = 8'h47 == _T_1[7:0] ? 8'h0 : _GEN_510; // @[Cat.scala 29:58]
  wire [7:0] _GEN_512 = 8'h48 == _T_1[7:0] ? 8'h0 : _GEN_511; // @[Cat.scala 29:58]
  wire [7:0] _GEN_513 = 8'h49 == _T_1[7:0] ? 8'h0 : _GEN_512; // @[Cat.scala 29:58]
  wire [7:0] _GEN_514 = 8'h4a == _T_1[7:0] ? 8'h0 : _GEN_513; // @[Cat.scala 29:58]
  wire [7:0] _GEN_515 = 8'h4b == _T_1[7:0] ? 8'h0 : _GEN_514; // @[Cat.scala 29:58]
  wire [7:0] _GEN_516 = 8'h4c == _T_1[7:0] ? 8'h0 : _GEN_515; // @[Cat.scala 29:58]
  wire [7:0] _GEN_517 = 8'h4d == _T_1[7:0] ? 8'h0 : _GEN_516; // @[Cat.scala 29:58]
  wire [7:0] _GEN_518 = 8'h4e == _T_1[7:0] ? 8'h0 : _GEN_517; // @[Cat.scala 29:58]
  wire [7:0] _GEN_519 = 8'h4f == _T_1[7:0] ? 8'h0 : _GEN_518; // @[Cat.scala 29:58]
  wire [7:0] _GEN_520 = 8'h50 == _T_1[7:0] ? 8'h0 : _GEN_519; // @[Cat.scala 29:58]
  wire [7:0] _GEN_521 = 8'h51 == _T_1[7:0] ? 8'h0 : _GEN_520; // @[Cat.scala 29:58]
  wire [7:0] _GEN_522 = 8'h52 == _T_1[7:0] ? 8'h0 : _GEN_521; // @[Cat.scala 29:58]
  wire [7:0] _GEN_523 = 8'h53 == _T_1[7:0] ? 8'h0 : _GEN_522; // @[Cat.scala 29:58]
  wire [7:0] _GEN_524 = 8'h54 == _T_1[7:0] ? 8'h0 : _GEN_523; // @[Cat.scala 29:58]
  wire [7:0] _GEN_525 = 8'h55 == _T_1[7:0] ? 8'h0 : _GEN_524; // @[Cat.scala 29:58]
  wire [7:0] _GEN_526 = 8'h56 == _T_1[7:0] ? 8'h0 : _GEN_525; // @[Cat.scala 29:58]
  wire [7:0] _GEN_527 = 8'h57 == _T_1[7:0] ? 8'h0 : _GEN_526; // @[Cat.scala 29:58]
  wire [7:0] _GEN_528 = 8'h58 == _T_1[7:0] ? 8'h0 : _GEN_527; // @[Cat.scala 29:58]
  wire [7:0] _GEN_529 = 8'h59 == _T_1[7:0] ? 8'h0 : _GEN_528; // @[Cat.scala 29:58]
  wire [7:0] _GEN_530 = 8'h5a == _T_1[7:0] ? 8'h0 : _GEN_529; // @[Cat.scala 29:58]
  wire [7:0] _GEN_531 = 8'h5b == _T_1[7:0] ? 8'h0 : _GEN_530; // @[Cat.scala 29:58]
  wire [7:0] _GEN_532 = 8'h5c == _T_1[7:0] ? 8'h0 : _GEN_531; // @[Cat.scala 29:58]
  wire [7:0] _GEN_533 = 8'h5d == _T_1[7:0] ? 8'h0 : _GEN_532; // @[Cat.scala 29:58]
  wire [7:0] _GEN_534 = 8'h5e == _T_1[7:0] ? 8'h0 : _GEN_533; // @[Cat.scala 29:58]
  wire [7:0] _GEN_535 = 8'h5f == _T_1[7:0] ? 8'h0 : _GEN_534; // @[Cat.scala 29:58]
  wire [7:0] _GEN_536 = 8'h60 == _T_1[7:0] ? 8'h0 : _GEN_535; // @[Cat.scala 29:58]
  wire [7:0] _GEN_537 = 8'h61 == _T_1[7:0] ? 8'h0 : _GEN_536; // @[Cat.scala 29:58]
  wire [7:0] _GEN_538 = 8'h62 == _T_1[7:0] ? 8'h0 : _GEN_537; // @[Cat.scala 29:58]
  wire [7:0] _GEN_539 = 8'h63 == _T_1[7:0] ? 8'h0 : _GEN_538; // @[Cat.scala 29:58]
  wire [7:0] _GEN_540 = 8'h64 == _T_1[7:0] ? 8'h0 : _GEN_539; // @[Cat.scala 29:58]
  wire [7:0] _GEN_541 = 8'h65 == _T_1[7:0] ? 8'h0 : _GEN_540; // @[Cat.scala 29:58]
  wire [7:0] _GEN_542 = 8'h66 == _T_1[7:0] ? 8'h0 : _GEN_541; // @[Cat.scala 29:58]
  wire [7:0] _GEN_543 = 8'h67 == _T_1[7:0] ? 8'h0 : _GEN_542; // @[Cat.scala 29:58]
  wire [7:0] _GEN_544 = 8'h68 == _T_1[7:0] ? 8'h0 : _GEN_543; // @[Cat.scala 29:58]
  wire [7:0] _GEN_545 = 8'h69 == _T_1[7:0] ? 8'h0 : _GEN_544; // @[Cat.scala 29:58]
  wire [7:0] _GEN_546 = 8'h6a == _T_1[7:0] ? 8'h0 : _GEN_545; // @[Cat.scala 29:58]
  wire [7:0] _GEN_547 = 8'h6b == _T_1[7:0] ? 8'h0 : _GEN_546; // @[Cat.scala 29:58]
  wire [7:0] _GEN_548 = 8'h6c == _T_1[7:0] ? 8'h0 : _GEN_547; // @[Cat.scala 29:58]
  wire [7:0] _GEN_549 = 8'h6d == _T_1[7:0] ? 8'h0 : _GEN_548; // @[Cat.scala 29:58]
  wire [7:0] _GEN_550 = 8'h6e == _T_1[7:0] ? 8'h0 : _GEN_549; // @[Cat.scala 29:58]
  wire [7:0] _GEN_551 = 8'h6f == _T_1[7:0] ? 8'h0 : _GEN_550; // @[Cat.scala 29:58]
  wire [7:0] _GEN_552 = 8'h70 == _T_1[7:0] ? 8'h0 : _GEN_551; // @[Cat.scala 29:58]
  wire [7:0] _GEN_553 = 8'h71 == _T_1[7:0] ? 8'h0 : _GEN_552; // @[Cat.scala 29:58]
  wire [7:0] _GEN_554 = 8'h72 == _T_1[7:0] ? 8'h0 : _GEN_553; // @[Cat.scala 29:58]
  wire [7:0] _GEN_555 = 8'h73 == _T_1[7:0] ? 8'h0 : _GEN_554; // @[Cat.scala 29:58]
  wire [7:0] _GEN_556 = 8'h74 == _T_1[7:0] ? 8'h0 : _GEN_555; // @[Cat.scala 29:58]
  wire [7:0] _GEN_557 = 8'h75 == _T_1[7:0] ? 8'h0 : _GEN_556; // @[Cat.scala 29:58]
  wire [7:0] _GEN_558 = 8'h76 == _T_1[7:0] ? 8'h0 : _GEN_557; // @[Cat.scala 29:58]
  wire [7:0] _GEN_559 = 8'h77 == _T_1[7:0] ? 8'h0 : _GEN_558; // @[Cat.scala 29:58]
  wire [7:0] _GEN_560 = 8'h78 == _T_1[7:0] ? 8'h0 : _GEN_559; // @[Cat.scala 29:58]
  wire [7:0] _GEN_561 = 8'h79 == _T_1[7:0] ? 8'h0 : _GEN_560; // @[Cat.scala 29:58]
  wire [7:0] _GEN_562 = 8'h7a == _T_1[7:0] ? 8'h0 : _GEN_561; // @[Cat.scala 29:58]
  wire [7:0] _GEN_563 = 8'h7b == _T_1[7:0] ? 8'h0 : _GEN_562; // @[Cat.scala 29:58]
  wire [7:0] _GEN_564 = 8'h7c == _T_1[7:0] ? 8'h0 : _GEN_563; // @[Cat.scala 29:58]
  wire [7:0] _GEN_565 = 8'h7d == _T_1[7:0] ? 8'h0 : _GEN_564; // @[Cat.scala 29:58]
  wire [7:0] _GEN_566 = 8'h7e == _T_1[7:0] ? 8'h0 : _GEN_565; // @[Cat.scala 29:58]
  wire [7:0] _GEN_567 = 8'h7f == _T_1[7:0] ? 8'h0 : _GEN_566; // @[Cat.scala 29:58]
  wire [7:0] _GEN_568 = 8'h80 == _T_1[7:0] ? 8'h0 : _GEN_567; // @[Cat.scala 29:58]
  wire [7:0] _GEN_569 = 8'h81 == _T_1[7:0] ? 8'h0 : _GEN_568; // @[Cat.scala 29:58]
  wire [7:0] _GEN_570 = 8'h82 == _T_1[7:0] ? 8'h0 : _GEN_569; // @[Cat.scala 29:58]
  wire [7:0] _GEN_571 = 8'h83 == _T_1[7:0] ? 8'h0 : _GEN_570; // @[Cat.scala 29:58]
  wire [7:0] _GEN_572 = 8'h84 == _T_1[7:0] ? 8'h0 : _GEN_571; // @[Cat.scala 29:58]
  wire [7:0] _GEN_573 = 8'h85 == _T_1[7:0] ? 8'h0 : _GEN_572; // @[Cat.scala 29:58]
  wire [7:0] _GEN_574 = 8'h86 == _T_1[7:0] ? 8'h0 : _GEN_573; // @[Cat.scala 29:58]
  wire [7:0] _GEN_575 = 8'h87 == _T_1[7:0] ? 8'h0 : _GEN_574; // @[Cat.scala 29:58]
  wire [7:0] _GEN_576 = 8'h88 == _T_1[7:0] ? 8'h0 : _GEN_575; // @[Cat.scala 29:58]
  wire [7:0] _GEN_577 = 8'h89 == _T_1[7:0] ? 8'h0 : _GEN_576; // @[Cat.scala 29:58]
  wire [7:0] _GEN_578 = 8'h8a == _T_1[7:0] ? 8'h0 : _GEN_577; // @[Cat.scala 29:58]
  wire [7:0] _GEN_579 = 8'h8b == _T_1[7:0] ? 8'h0 : _GEN_578; // @[Cat.scala 29:58]
  wire [7:0] _GEN_580 = 8'h8c == _T_1[7:0] ? 8'h0 : _GEN_579; // @[Cat.scala 29:58]
  wire [7:0] _GEN_581 = 8'h8d == _T_1[7:0] ? 8'h0 : _GEN_580; // @[Cat.scala 29:58]
  wire [7:0] _GEN_582 = 8'h8e == _T_1[7:0] ? 8'h0 : _GEN_581; // @[Cat.scala 29:58]
  wire [7:0] _GEN_583 = 8'h8f == _T_1[7:0] ? 8'h0 : _GEN_582; // @[Cat.scala 29:58]
  wire [7:0] _GEN_584 = 8'h90 == _T_1[7:0] ? 8'h0 : _GEN_583; // @[Cat.scala 29:58]
  wire [7:0] _GEN_585 = 8'h91 == _T_1[7:0] ? 8'h0 : _GEN_584; // @[Cat.scala 29:58]
  wire [7:0] _GEN_586 = 8'h92 == _T_1[7:0] ? 8'h0 : _GEN_585; // @[Cat.scala 29:58]
  wire [7:0] _GEN_587 = 8'h93 == _T_1[7:0] ? 8'h0 : _GEN_586; // @[Cat.scala 29:58]
  wire [7:0] _GEN_588 = 8'h94 == _T_1[7:0] ? 8'h0 : _GEN_587; // @[Cat.scala 29:58]
  wire [7:0] _GEN_589 = 8'h95 == _T_1[7:0] ? 8'h0 : _GEN_588; // @[Cat.scala 29:58]
  wire [7:0] _GEN_590 = 8'h96 == _T_1[7:0] ? 8'h0 : _GEN_589; // @[Cat.scala 29:58]
  wire [7:0] _GEN_591 = 8'h97 == _T_1[7:0] ? 8'h0 : _GEN_590; // @[Cat.scala 29:58]
  wire [7:0] _GEN_592 = 8'h98 == _T_1[7:0] ? 8'h0 : _GEN_591; // @[Cat.scala 29:58]
  wire [7:0] _GEN_593 = 8'h99 == _T_1[7:0] ? 8'h0 : _GEN_592; // @[Cat.scala 29:58]
  wire [7:0] _GEN_594 = 8'h9a == _T_1[7:0] ? 8'h0 : _GEN_593; // @[Cat.scala 29:58]
  wire [7:0] _GEN_595 = 8'h9b == _T_1[7:0] ? 8'h0 : _GEN_594; // @[Cat.scala 29:58]
  wire [7:0] _GEN_596 = 8'h9c == _T_1[7:0] ? 8'h0 : _GEN_595; // @[Cat.scala 29:58]
  wire [7:0] _GEN_597 = 8'h9d == _T_1[7:0] ? 8'h0 : _GEN_596; // @[Cat.scala 29:58]
  wire [7:0] _GEN_598 = 8'h9e == _T_1[7:0] ? 8'h0 : _GEN_597; // @[Cat.scala 29:58]
  wire [7:0] _GEN_599 = 8'h9f == _T_1[7:0] ? 8'h0 : _GEN_598; // @[Cat.scala 29:58]
  wire [7:0] _GEN_600 = 8'ha0 == _T_1[7:0] ? 8'h0 : _GEN_599; // @[Cat.scala 29:58]
  wire [7:0] _GEN_601 = 8'ha1 == _T_1[7:0] ? 8'h0 : _GEN_600; // @[Cat.scala 29:58]
  wire [7:0] _GEN_602 = 8'ha2 == _T_1[7:0] ? 8'h0 : _GEN_601; // @[Cat.scala 29:58]
  wire [7:0] _GEN_603 = 8'ha3 == _T_1[7:0] ? 8'h0 : _GEN_602; // @[Cat.scala 29:58]
  wire [7:0] _GEN_604 = 8'ha4 == _T_1[7:0] ? 8'h0 : _GEN_603; // @[Cat.scala 29:58]
  wire [7:0] _GEN_605 = 8'ha5 == _T_1[7:0] ? 8'h0 : _GEN_604; // @[Cat.scala 29:58]
  wire [7:0] _GEN_606 = 8'ha6 == _T_1[7:0] ? 8'h0 : _GEN_605; // @[Cat.scala 29:58]
  wire [7:0] _GEN_607 = 8'ha7 == _T_1[7:0] ? 8'h0 : _GEN_606; // @[Cat.scala 29:58]
  wire [7:0] _GEN_608 = 8'ha8 == _T_1[7:0] ? 8'h0 : _GEN_607; // @[Cat.scala 29:58]
  wire [7:0] _GEN_609 = 8'ha9 == _T_1[7:0] ? 8'h0 : _GEN_608; // @[Cat.scala 29:58]
  wire [7:0] _GEN_610 = 8'haa == _T_1[7:0] ? 8'h0 : _GEN_609; // @[Cat.scala 29:58]
  wire [7:0] _GEN_611 = 8'hab == _T_1[7:0] ? 8'h0 : _GEN_610; // @[Cat.scala 29:58]
  wire [7:0] _GEN_612 = 8'hac == _T_1[7:0] ? 8'h0 : _GEN_611; // @[Cat.scala 29:58]
  wire [7:0] _GEN_613 = 8'had == _T_1[7:0] ? 8'h0 : _GEN_612; // @[Cat.scala 29:58]
  wire [7:0] _GEN_614 = 8'hae == _T_1[7:0] ? 8'h0 : _GEN_613; // @[Cat.scala 29:58]
  wire [7:0] _GEN_615 = 8'haf == _T_1[7:0] ? 8'h0 : _GEN_614; // @[Cat.scala 29:58]
  wire [7:0] _GEN_616 = 8'hb0 == _T_1[7:0] ? 8'h0 : _GEN_615; // @[Cat.scala 29:58]
  wire [7:0] _GEN_617 = 8'hb1 == _T_1[7:0] ? 8'h0 : _GEN_616; // @[Cat.scala 29:58]
  wire [7:0] _GEN_618 = 8'hb2 == _T_1[7:0] ? 8'h0 : _GEN_617; // @[Cat.scala 29:58]
  wire [7:0] _GEN_619 = 8'hb3 == _T_1[7:0] ? 8'h0 : _GEN_618; // @[Cat.scala 29:58]
  wire [7:0] _GEN_620 = 8'hb4 == _T_1[7:0] ? 8'h0 : _GEN_619; // @[Cat.scala 29:58]
  wire [7:0] _GEN_621 = 8'hb5 == _T_1[7:0] ? 8'h0 : _GEN_620; // @[Cat.scala 29:58]
  wire [7:0] _GEN_622 = 8'hb6 == _T_1[7:0] ? 8'h0 : _GEN_621; // @[Cat.scala 29:58]
  wire [7:0] _GEN_623 = 8'hb7 == _T_1[7:0] ? 8'h0 : _GEN_622; // @[Cat.scala 29:58]
  wire [7:0] _GEN_624 = 8'hb8 == _T_1[7:0] ? 8'h0 : _GEN_623; // @[Cat.scala 29:58]
  wire [7:0] _GEN_625 = 8'hb9 == _T_1[7:0] ? 8'h0 : _GEN_624; // @[Cat.scala 29:58]
  wire [7:0] _GEN_626 = 8'hba == _T_1[7:0] ? 8'h0 : _GEN_625; // @[Cat.scala 29:58]
  wire [7:0] _GEN_627 = 8'hbb == _T_1[7:0] ? 8'h0 : _GEN_626; // @[Cat.scala 29:58]
  wire [7:0] _GEN_628 = 8'hbc == _T_1[7:0] ? 8'h0 : _GEN_627; // @[Cat.scala 29:58]
  wire [7:0] _GEN_629 = 8'hbd == _T_1[7:0] ? 8'h0 : _GEN_628; // @[Cat.scala 29:58]
  wire [7:0] _GEN_630 = 8'hbe == _T_1[7:0] ? 8'h0 : _GEN_629; // @[Cat.scala 29:58]
  wire [7:0] _GEN_631 = 8'hbf == _T_1[7:0] ? 8'h0 : _GEN_630; // @[Cat.scala 29:58]
  wire [7:0] _GEN_632 = 8'hc0 == _T_1[7:0] ? 8'h0 : _GEN_631; // @[Cat.scala 29:58]
  wire [7:0] _GEN_633 = 8'hc1 == _T_1[7:0] ? 8'h0 : _GEN_632; // @[Cat.scala 29:58]
  wire [7:0] _GEN_634 = 8'hc2 == _T_1[7:0] ? 8'h0 : _GEN_633; // @[Cat.scala 29:58]
  wire [7:0] _GEN_635 = 8'hc3 == _T_1[7:0] ? 8'h0 : _GEN_634; // @[Cat.scala 29:58]
  wire [7:0] _GEN_636 = 8'hc4 == _T_1[7:0] ? 8'h0 : _GEN_635; // @[Cat.scala 29:58]
  wire [7:0] _GEN_637 = 8'hc5 == _T_1[7:0] ? 8'h0 : _GEN_636; // @[Cat.scala 29:58]
  wire [7:0] _GEN_638 = 8'hc6 == _T_1[7:0] ? 8'h0 : _GEN_637; // @[Cat.scala 29:58]
  wire [7:0] _GEN_639 = 8'hc7 == _T_1[7:0] ? 8'h0 : _GEN_638; // @[Cat.scala 29:58]
  wire [7:0] _GEN_640 = 8'hc8 == _T_1[7:0] ? 8'h0 : _GEN_639; // @[Cat.scala 29:58]
  wire [7:0] _GEN_641 = 8'hc9 == _T_1[7:0] ? 8'h0 : _GEN_640; // @[Cat.scala 29:58]
  wire [7:0] _GEN_642 = 8'hca == _T_1[7:0] ? 8'h0 : _GEN_641; // @[Cat.scala 29:58]
  wire [7:0] _GEN_643 = 8'hcb == _T_1[7:0] ? 8'h0 : _GEN_642; // @[Cat.scala 29:58]
  wire [7:0] _GEN_644 = 8'hcc == _T_1[7:0] ? 8'h0 : _GEN_643; // @[Cat.scala 29:58]
  wire [7:0] _GEN_645 = 8'hcd == _T_1[7:0] ? 8'h0 : _GEN_644; // @[Cat.scala 29:58]
  wire [7:0] _GEN_646 = 8'hce == _T_1[7:0] ? 8'h0 : _GEN_645; // @[Cat.scala 29:58]
  wire [7:0] _GEN_647 = 8'hcf == _T_1[7:0] ? 8'h0 : _GEN_646; // @[Cat.scala 29:58]
  wire [7:0] _GEN_648 = 8'hd0 == _T_1[7:0] ? 8'h0 : _GEN_647; // @[Cat.scala 29:58]
  wire [7:0] _GEN_649 = 8'hd1 == _T_1[7:0] ? 8'h0 : _GEN_648; // @[Cat.scala 29:58]
  wire [7:0] _GEN_650 = 8'hd2 == _T_1[7:0] ? 8'h0 : _GEN_649; // @[Cat.scala 29:58]
  wire [7:0] _GEN_651 = 8'hd3 == _T_1[7:0] ? 8'h0 : _GEN_650; // @[Cat.scala 29:58]
  wire [7:0] _GEN_652 = 8'hd4 == _T_1[7:0] ? 8'h0 : _GEN_651; // @[Cat.scala 29:58]
  wire [7:0] _GEN_653 = 8'hd5 == _T_1[7:0] ? 8'h0 : _GEN_652; // @[Cat.scala 29:58]
  wire [7:0] _GEN_654 = 8'hd6 == _T_1[7:0] ? 8'h0 : _GEN_653; // @[Cat.scala 29:58]
  wire [7:0] _GEN_655 = 8'hd7 == _T_1[7:0] ? 8'h0 : _GEN_654; // @[Cat.scala 29:58]
  wire [7:0] _GEN_656 = 8'hd8 == _T_1[7:0] ? 8'h0 : _GEN_655; // @[Cat.scala 29:58]
  wire [7:0] _GEN_657 = 8'hd9 == _T_1[7:0] ? 8'h0 : _GEN_656; // @[Cat.scala 29:58]
  wire [7:0] _GEN_658 = 8'hda == _T_1[7:0] ? 8'h0 : _GEN_657; // @[Cat.scala 29:58]
  wire [7:0] _GEN_659 = 8'hdb == _T_1[7:0] ? 8'h0 : _GEN_658; // @[Cat.scala 29:58]
  wire [7:0] _GEN_661 = 8'h1 == _T_4[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_662 = 8'h2 == _T_4[7:0] ? 8'h0 : _GEN_661; // @[Cat.scala 29:58]
  wire [7:0] _GEN_663 = 8'h3 == _T_4[7:0] ? 8'hfe : _GEN_662; // @[Cat.scala 29:58]
  wire [7:0] _GEN_664 = 8'h4 == _T_4[7:0] ? 8'h93 : _GEN_663; // @[Cat.scala 29:58]
  wire [7:0] _GEN_665 = 8'h5 == _T_4[7:0] ? 8'h5 : _GEN_664; // @[Cat.scala 29:58]
  wire [7:0] _GEN_666 = 8'h6 == _T_4[7:0] ? 8'h0 : _GEN_665; // @[Cat.scala 29:58]
  wire [7:0] _GEN_667 = 8'h7 == _T_4[7:0] ? 8'hfc : _GEN_666; // @[Cat.scala 29:58]
  wire [7:0] _GEN_668 = 8'h8 == _T_4[7:0] ? 8'h33 : _GEN_667; // @[Cat.scala 29:58]
  wire [7:0] _GEN_669 = 8'h9 == _T_4[7:0] ? 8'h6 : _GEN_668; // @[Cat.scala 29:58]
  wire [7:0] _GEN_670 = 8'ha == _T_4[7:0] ? 8'hb5 : _GEN_669; // @[Cat.scala 29:58]
  wire [7:0] _GEN_671 = 8'hb == _T_4[7:0] ? 8'h0 : _GEN_670; // @[Cat.scala 29:58]
  wire [7:0] _GEN_672 = 8'hc == _T_4[7:0] ? 8'h13 : _GEN_671; // @[Cat.scala 29:58]
  wire [7:0] _GEN_673 = 8'hd == _T_4[7:0] ? 8'h5 : _GEN_672; // @[Cat.scala 29:58]
  wire [7:0] _GEN_674 = 8'he == _T_4[7:0] ? 8'ha0 : _GEN_673; // @[Cat.scala 29:58]
  wire [7:0] _GEN_675 = 8'hf == _T_4[7:0] ? 8'h0 : _GEN_674; // @[Cat.scala 29:58]
  wire [7:0] _GEN_676 = 8'h10 == _T_4[7:0] ? 8'h73 : _GEN_675; // @[Cat.scala 29:58]
  wire [7:0] _GEN_677 = 8'h11 == _T_4[7:0] ? 8'h0 : _GEN_676; // @[Cat.scala 29:58]
  wire [7:0] _GEN_678 = 8'h12 == _T_4[7:0] ? 8'h0 : _GEN_677; // @[Cat.scala 29:58]
  wire [7:0] _GEN_679 = 8'h13 == _T_4[7:0] ? 8'h0 : _GEN_678; // @[Cat.scala 29:58]
  wire [7:0] _GEN_680 = 8'h14 == _T_4[7:0] ? 8'h0 : _GEN_679; // @[Cat.scala 29:58]
  wire [7:0] _GEN_681 = 8'h15 == _T_4[7:0] ? 8'h0 : _GEN_680; // @[Cat.scala 29:58]
  wire [7:0] _GEN_682 = 8'h16 == _T_4[7:0] ? 8'h0 : _GEN_681; // @[Cat.scala 29:58]
  wire [7:0] _GEN_683 = 8'h17 == _T_4[7:0] ? 8'h0 : _GEN_682; // @[Cat.scala 29:58]
  wire [7:0] _GEN_684 = 8'h18 == _T_4[7:0] ? 8'h0 : _GEN_683; // @[Cat.scala 29:58]
  wire [7:0] _GEN_685 = 8'h19 == _T_4[7:0] ? 8'h0 : _GEN_684; // @[Cat.scala 29:58]
  wire [7:0] _GEN_686 = 8'h1a == _T_4[7:0] ? 8'h0 : _GEN_685; // @[Cat.scala 29:58]
  wire [7:0] _GEN_687 = 8'h1b == _T_4[7:0] ? 8'h0 : _GEN_686; // @[Cat.scala 29:58]
  wire [7:0] _GEN_688 = 8'h1c == _T_4[7:0] ? 8'h0 : _GEN_687; // @[Cat.scala 29:58]
  wire [7:0] _GEN_689 = 8'h1d == _T_4[7:0] ? 8'h0 : _GEN_688; // @[Cat.scala 29:58]
  wire [7:0] _GEN_690 = 8'h1e == _T_4[7:0] ? 8'h0 : _GEN_689; // @[Cat.scala 29:58]
  wire [7:0] _GEN_691 = 8'h1f == _T_4[7:0] ? 8'h0 : _GEN_690; // @[Cat.scala 29:58]
  wire [7:0] _GEN_692 = 8'h20 == _T_4[7:0] ? 8'h0 : _GEN_691; // @[Cat.scala 29:58]
  wire [7:0] _GEN_693 = 8'h21 == _T_4[7:0] ? 8'h0 : _GEN_692; // @[Cat.scala 29:58]
  wire [7:0] _GEN_694 = 8'h22 == _T_4[7:0] ? 8'h0 : _GEN_693; // @[Cat.scala 29:58]
  wire [7:0] _GEN_695 = 8'h23 == _T_4[7:0] ? 8'h0 : _GEN_694; // @[Cat.scala 29:58]
  wire [7:0] _GEN_696 = 8'h24 == _T_4[7:0] ? 8'h0 : _GEN_695; // @[Cat.scala 29:58]
  wire [7:0] _GEN_697 = 8'h25 == _T_4[7:0] ? 8'h0 : _GEN_696; // @[Cat.scala 29:58]
  wire [7:0] _GEN_698 = 8'h26 == _T_4[7:0] ? 8'h0 : _GEN_697; // @[Cat.scala 29:58]
  wire [7:0] _GEN_699 = 8'h27 == _T_4[7:0] ? 8'h0 : _GEN_698; // @[Cat.scala 29:58]
  wire [7:0] _GEN_700 = 8'h28 == _T_4[7:0] ? 8'h0 : _GEN_699; // @[Cat.scala 29:58]
  wire [7:0] _GEN_701 = 8'h29 == _T_4[7:0] ? 8'h0 : _GEN_700; // @[Cat.scala 29:58]
  wire [7:0] _GEN_702 = 8'h2a == _T_4[7:0] ? 8'h0 : _GEN_701; // @[Cat.scala 29:58]
  wire [7:0] _GEN_703 = 8'h2b == _T_4[7:0] ? 8'h0 : _GEN_702; // @[Cat.scala 29:58]
  wire [7:0] _GEN_704 = 8'h2c == _T_4[7:0] ? 8'h0 : _GEN_703; // @[Cat.scala 29:58]
  wire [7:0] _GEN_705 = 8'h2d == _T_4[7:0] ? 8'h0 : _GEN_704; // @[Cat.scala 29:58]
  wire [7:0] _GEN_706 = 8'h2e == _T_4[7:0] ? 8'h0 : _GEN_705; // @[Cat.scala 29:58]
  wire [7:0] _GEN_707 = 8'h2f == _T_4[7:0] ? 8'h0 : _GEN_706; // @[Cat.scala 29:58]
  wire [7:0] _GEN_708 = 8'h30 == _T_4[7:0] ? 8'h0 : _GEN_707; // @[Cat.scala 29:58]
  wire [7:0] _GEN_709 = 8'h31 == _T_4[7:0] ? 8'h0 : _GEN_708; // @[Cat.scala 29:58]
  wire [7:0] _GEN_710 = 8'h32 == _T_4[7:0] ? 8'h0 : _GEN_709; // @[Cat.scala 29:58]
  wire [7:0] _GEN_711 = 8'h33 == _T_4[7:0] ? 8'h0 : _GEN_710; // @[Cat.scala 29:58]
  wire [7:0] _GEN_712 = 8'h34 == _T_4[7:0] ? 8'h0 : _GEN_711; // @[Cat.scala 29:58]
  wire [7:0] _GEN_713 = 8'h35 == _T_4[7:0] ? 8'h0 : _GEN_712; // @[Cat.scala 29:58]
  wire [7:0] _GEN_714 = 8'h36 == _T_4[7:0] ? 8'h0 : _GEN_713; // @[Cat.scala 29:58]
  wire [7:0] _GEN_715 = 8'h37 == _T_4[7:0] ? 8'h0 : _GEN_714; // @[Cat.scala 29:58]
  wire [7:0] _GEN_716 = 8'h38 == _T_4[7:0] ? 8'h0 : _GEN_715; // @[Cat.scala 29:58]
  wire [7:0] _GEN_717 = 8'h39 == _T_4[7:0] ? 8'h0 : _GEN_716; // @[Cat.scala 29:58]
  wire [7:0] _GEN_718 = 8'h3a == _T_4[7:0] ? 8'h0 : _GEN_717; // @[Cat.scala 29:58]
  wire [7:0] _GEN_719 = 8'h3b == _T_4[7:0] ? 8'h0 : _GEN_718; // @[Cat.scala 29:58]
  wire [7:0] _GEN_720 = 8'h3c == _T_4[7:0] ? 8'h0 : _GEN_719; // @[Cat.scala 29:58]
  wire [7:0] _GEN_721 = 8'h3d == _T_4[7:0] ? 8'h0 : _GEN_720; // @[Cat.scala 29:58]
  wire [7:0] _GEN_722 = 8'h3e == _T_4[7:0] ? 8'h0 : _GEN_721; // @[Cat.scala 29:58]
  wire [7:0] _GEN_723 = 8'h3f == _T_4[7:0] ? 8'h0 : _GEN_722; // @[Cat.scala 29:58]
  wire [7:0] _GEN_724 = 8'h40 == _T_4[7:0] ? 8'h0 : _GEN_723; // @[Cat.scala 29:58]
  wire [7:0] _GEN_725 = 8'h41 == _T_4[7:0] ? 8'h0 : _GEN_724; // @[Cat.scala 29:58]
  wire [7:0] _GEN_726 = 8'h42 == _T_4[7:0] ? 8'h0 : _GEN_725; // @[Cat.scala 29:58]
  wire [7:0] _GEN_727 = 8'h43 == _T_4[7:0] ? 8'h0 : _GEN_726; // @[Cat.scala 29:58]
  wire [7:0] _GEN_728 = 8'h44 == _T_4[7:0] ? 8'h0 : _GEN_727; // @[Cat.scala 29:58]
  wire [7:0] _GEN_729 = 8'h45 == _T_4[7:0] ? 8'h0 : _GEN_728; // @[Cat.scala 29:58]
  wire [7:0] _GEN_730 = 8'h46 == _T_4[7:0] ? 8'h0 : _GEN_729; // @[Cat.scala 29:58]
  wire [7:0] _GEN_731 = 8'h47 == _T_4[7:0] ? 8'h0 : _GEN_730; // @[Cat.scala 29:58]
  wire [7:0] _GEN_732 = 8'h48 == _T_4[7:0] ? 8'h0 : _GEN_731; // @[Cat.scala 29:58]
  wire [7:0] _GEN_733 = 8'h49 == _T_4[7:0] ? 8'h0 : _GEN_732; // @[Cat.scala 29:58]
  wire [7:0] _GEN_734 = 8'h4a == _T_4[7:0] ? 8'h0 : _GEN_733; // @[Cat.scala 29:58]
  wire [7:0] _GEN_735 = 8'h4b == _T_4[7:0] ? 8'h0 : _GEN_734; // @[Cat.scala 29:58]
  wire [7:0] _GEN_736 = 8'h4c == _T_4[7:0] ? 8'h0 : _GEN_735; // @[Cat.scala 29:58]
  wire [7:0] _GEN_737 = 8'h4d == _T_4[7:0] ? 8'h0 : _GEN_736; // @[Cat.scala 29:58]
  wire [7:0] _GEN_738 = 8'h4e == _T_4[7:0] ? 8'h0 : _GEN_737; // @[Cat.scala 29:58]
  wire [7:0] _GEN_739 = 8'h4f == _T_4[7:0] ? 8'h0 : _GEN_738; // @[Cat.scala 29:58]
  wire [7:0] _GEN_740 = 8'h50 == _T_4[7:0] ? 8'h0 : _GEN_739; // @[Cat.scala 29:58]
  wire [7:0] _GEN_741 = 8'h51 == _T_4[7:0] ? 8'h0 : _GEN_740; // @[Cat.scala 29:58]
  wire [7:0] _GEN_742 = 8'h52 == _T_4[7:0] ? 8'h0 : _GEN_741; // @[Cat.scala 29:58]
  wire [7:0] _GEN_743 = 8'h53 == _T_4[7:0] ? 8'h0 : _GEN_742; // @[Cat.scala 29:58]
  wire [7:0] _GEN_744 = 8'h54 == _T_4[7:0] ? 8'h0 : _GEN_743; // @[Cat.scala 29:58]
  wire [7:0] _GEN_745 = 8'h55 == _T_4[7:0] ? 8'h0 : _GEN_744; // @[Cat.scala 29:58]
  wire [7:0] _GEN_746 = 8'h56 == _T_4[7:0] ? 8'h0 : _GEN_745; // @[Cat.scala 29:58]
  wire [7:0] _GEN_747 = 8'h57 == _T_4[7:0] ? 8'h0 : _GEN_746; // @[Cat.scala 29:58]
  wire [7:0] _GEN_748 = 8'h58 == _T_4[7:0] ? 8'h0 : _GEN_747; // @[Cat.scala 29:58]
  wire [7:0] _GEN_749 = 8'h59 == _T_4[7:0] ? 8'h0 : _GEN_748; // @[Cat.scala 29:58]
  wire [7:0] _GEN_750 = 8'h5a == _T_4[7:0] ? 8'h0 : _GEN_749; // @[Cat.scala 29:58]
  wire [7:0] _GEN_751 = 8'h5b == _T_4[7:0] ? 8'h0 : _GEN_750; // @[Cat.scala 29:58]
  wire [7:0] _GEN_752 = 8'h5c == _T_4[7:0] ? 8'h0 : _GEN_751; // @[Cat.scala 29:58]
  wire [7:0] _GEN_753 = 8'h5d == _T_4[7:0] ? 8'h0 : _GEN_752; // @[Cat.scala 29:58]
  wire [7:0] _GEN_754 = 8'h5e == _T_4[7:0] ? 8'h0 : _GEN_753; // @[Cat.scala 29:58]
  wire [7:0] _GEN_755 = 8'h5f == _T_4[7:0] ? 8'h0 : _GEN_754; // @[Cat.scala 29:58]
  wire [7:0] _GEN_756 = 8'h60 == _T_4[7:0] ? 8'h0 : _GEN_755; // @[Cat.scala 29:58]
  wire [7:0] _GEN_757 = 8'h61 == _T_4[7:0] ? 8'h0 : _GEN_756; // @[Cat.scala 29:58]
  wire [7:0] _GEN_758 = 8'h62 == _T_4[7:0] ? 8'h0 : _GEN_757; // @[Cat.scala 29:58]
  wire [7:0] _GEN_759 = 8'h63 == _T_4[7:0] ? 8'h0 : _GEN_758; // @[Cat.scala 29:58]
  wire [7:0] _GEN_760 = 8'h64 == _T_4[7:0] ? 8'h0 : _GEN_759; // @[Cat.scala 29:58]
  wire [7:0] _GEN_761 = 8'h65 == _T_4[7:0] ? 8'h0 : _GEN_760; // @[Cat.scala 29:58]
  wire [7:0] _GEN_762 = 8'h66 == _T_4[7:0] ? 8'h0 : _GEN_761; // @[Cat.scala 29:58]
  wire [7:0] _GEN_763 = 8'h67 == _T_4[7:0] ? 8'h0 : _GEN_762; // @[Cat.scala 29:58]
  wire [7:0] _GEN_764 = 8'h68 == _T_4[7:0] ? 8'h0 : _GEN_763; // @[Cat.scala 29:58]
  wire [7:0] _GEN_765 = 8'h69 == _T_4[7:0] ? 8'h0 : _GEN_764; // @[Cat.scala 29:58]
  wire [7:0] _GEN_766 = 8'h6a == _T_4[7:0] ? 8'h0 : _GEN_765; // @[Cat.scala 29:58]
  wire [7:0] _GEN_767 = 8'h6b == _T_4[7:0] ? 8'h0 : _GEN_766; // @[Cat.scala 29:58]
  wire [7:0] _GEN_768 = 8'h6c == _T_4[7:0] ? 8'h0 : _GEN_767; // @[Cat.scala 29:58]
  wire [7:0] _GEN_769 = 8'h6d == _T_4[7:0] ? 8'h0 : _GEN_768; // @[Cat.scala 29:58]
  wire [7:0] _GEN_770 = 8'h6e == _T_4[7:0] ? 8'h0 : _GEN_769; // @[Cat.scala 29:58]
  wire [7:0] _GEN_771 = 8'h6f == _T_4[7:0] ? 8'h0 : _GEN_770; // @[Cat.scala 29:58]
  wire [7:0] _GEN_772 = 8'h70 == _T_4[7:0] ? 8'h0 : _GEN_771; // @[Cat.scala 29:58]
  wire [7:0] _GEN_773 = 8'h71 == _T_4[7:0] ? 8'h0 : _GEN_772; // @[Cat.scala 29:58]
  wire [7:0] _GEN_774 = 8'h72 == _T_4[7:0] ? 8'h0 : _GEN_773; // @[Cat.scala 29:58]
  wire [7:0] _GEN_775 = 8'h73 == _T_4[7:0] ? 8'h0 : _GEN_774; // @[Cat.scala 29:58]
  wire [7:0] _GEN_776 = 8'h74 == _T_4[7:0] ? 8'h0 : _GEN_775; // @[Cat.scala 29:58]
  wire [7:0] _GEN_777 = 8'h75 == _T_4[7:0] ? 8'h0 : _GEN_776; // @[Cat.scala 29:58]
  wire [7:0] _GEN_778 = 8'h76 == _T_4[7:0] ? 8'h0 : _GEN_777; // @[Cat.scala 29:58]
  wire [7:0] _GEN_779 = 8'h77 == _T_4[7:0] ? 8'h0 : _GEN_778; // @[Cat.scala 29:58]
  wire [7:0] _GEN_780 = 8'h78 == _T_4[7:0] ? 8'h0 : _GEN_779; // @[Cat.scala 29:58]
  wire [7:0] _GEN_781 = 8'h79 == _T_4[7:0] ? 8'h0 : _GEN_780; // @[Cat.scala 29:58]
  wire [7:0] _GEN_782 = 8'h7a == _T_4[7:0] ? 8'h0 : _GEN_781; // @[Cat.scala 29:58]
  wire [7:0] _GEN_783 = 8'h7b == _T_4[7:0] ? 8'h0 : _GEN_782; // @[Cat.scala 29:58]
  wire [7:0] _GEN_784 = 8'h7c == _T_4[7:0] ? 8'h0 : _GEN_783; // @[Cat.scala 29:58]
  wire [7:0] _GEN_785 = 8'h7d == _T_4[7:0] ? 8'h0 : _GEN_784; // @[Cat.scala 29:58]
  wire [7:0] _GEN_786 = 8'h7e == _T_4[7:0] ? 8'h0 : _GEN_785; // @[Cat.scala 29:58]
  wire [7:0] _GEN_787 = 8'h7f == _T_4[7:0] ? 8'h0 : _GEN_786; // @[Cat.scala 29:58]
  wire [7:0] _GEN_788 = 8'h80 == _T_4[7:0] ? 8'h0 : _GEN_787; // @[Cat.scala 29:58]
  wire [7:0] _GEN_789 = 8'h81 == _T_4[7:0] ? 8'h0 : _GEN_788; // @[Cat.scala 29:58]
  wire [7:0] _GEN_790 = 8'h82 == _T_4[7:0] ? 8'h0 : _GEN_789; // @[Cat.scala 29:58]
  wire [7:0] _GEN_791 = 8'h83 == _T_4[7:0] ? 8'h0 : _GEN_790; // @[Cat.scala 29:58]
  wire [7:0] _GEN_792 = 8'h84 == _T_4[7:0] ? 8'h0 : _GEN_791; // @[Cat.scala 29:58]
  wire [7:0] _GEN_793 = 8'h85 == _T_4[7:0] ? 8'h0 : _GEN_792; // @[Cat.scala 29:58]
  wire [7:0] _GEN_794 = 8'h86 == _T_4[7:0] ? 8'h0 : _GEN_793; // @[Cat.scala 29:58]
  wire [7:0] _GEN_795 = 8'h87 == _T_4[7:0] ? 8'h0 : _GEN_794; // @[Cat.scala 29:58]
  wire [7:0] _GEN_796 = 8'h88 == _T_4[7:0] ? 8'h0 : _GEN_795; // @[Cat.scala 29:58]
  wire [7:0] _GEN_797 = 8'h89 == _T_4[7:0] ? 8'h0 : _GEN_796; // @[Cat.scala 29:58]
  wire [7:0] _GEN_798 = 8'h8a == _T_4[7:0] ? 8'h0 : _GEN_797; // @[Cat.scala 29:58]
  wire [7:0] _GEN_799 = 8'h8b == _T_4[7:0] ? 8'h0 : _GEN_798; // @[Cat.scala 29:58]
  wire [7:0] _GEN_800 = 8'h8c == _T_4[7:0] ? 8'h0 : _GEN_799; // @[Cat.scala 29:58]
  wire [7:0] _GEN_801 = 8'h8d == _T_4[7:0] ? 8'h0 : _GEN_800; // @[Cat.scala 29:58]
  wire [7:0] _GEN_802 = 8'h8e == _T_4[7:0] ? 8'h0 : _GEN_801; // @[Cat.scala 29:58]
  wire [7:0] _GEN_803 = 8'h8f == _T_4[7:0] ? 8'h0 : _GEN_802; // @[Cat.scala 29:58]
  wire [7:0] _GEN_804 = 8'h90 == _T_4[7:0] ? 8'h0 : _GEN_803; // @[Cat.scala 29:58]
  wire [7:0] _GEN_805 = 8'h91 == _T_4[7:0] ? 8'h0 : _GEN_804; // @[Cat.scala 29:58]
  wire [7:0] _GEN_806 = 8'h92 == _T_4[7:0] ? 8'h0 : _GEN_805; // @[Cat.scala 29:58]
  wire [7:0] _GEN_807 = 8'h93 == _T_4[7:0] ? 8'h0 : _GEN_806; // @[Cat.scala 29:58]
  wire [7:0] _GEN_808 = 8'h94 == _T_4[7:0] ? 8'h0 : _GEN_807; // @[Cat.scala 29:58]
  wire [7:0] _GEN_809 = 8'h95 == _T_4[7:0] ? 8'h0 : _GEN_808; // @[Cat.scala 29:58]
  wire [7:0] _GEN_810 = 8'h96 == _T_4[7:0] ? 8'h0 : _GEN_809; // @[Cat.scala 29:58]
  wire [7:0] _GEN_811 = 8'h97 == _T_4[7:0] ? 8'h0 : _GEN_810; // @[Cat.scala 29:58]
  wire [7:0] _GEN_812 = 8'h98 == _T_4[7:0] ? 8'h0 : _GEN_811; // @[Cat.scala 29:58]
  wire [7:0] _GEN_813 = 8'h99 == _T_4[7:0] ? 8'h0 : _GEN_812; // @[Cat.scala 29:58]
  wire [7:0] _GEN_814 = 8'h9a == _T_4[7:0] ? 8'h0 : _GEN_813; // @[Cat.scala 29:58]
  wire [7:0] _GEN_815 = 8'h9b == _T_4[7:0] ? 8'h0 : _GEN_814; // @[Cat.scala 29:58]
  wire [7:0] _GEN_816 = 8'h9c == _T_4[7:0] ? 8'h0 : _GEN_815; // @[Cat.scala 29:58]
  wire [7:0] _GEN_817 = 8'h9d == _T_4[7:0] ? 8'h0 : _GEN_816; // @[Cat.scala 29:58]
  wire [7:0] _GEN_818 = 8'h9e == _T_4[7:0] ? 8'h0 : _GEN_817; // @[Cat.scala 29:58]
  wire [7:0] _GEN_819 = 8'h9f == _T_4[7:0] ? 8'h0 : _GEN_818; // @[Cat.scala 29:58]
  wire [7:0] _GEN_820 = 8'ha0 == _T_4[7:0] ? 8'h0 : _GEN_819; // @[Cat.scala 29:58]
  wire [7:0] _GEN_821 = 8'ha1 == _T_4[7:0] ? 8'h0 : _GEN_820; // @[Cat.scala 29:58]
  wire [7:0] _GEN_822 = 8'ha2 == _T_4[7:0] ? 8'h0 : _GEN_821; // @[Cat.scala 29:58]
  wire [7:0] _GEN_823 = 8'ha3 == _T_4[7:0] ? 8'h0 : _GEN_822; // @[Cat.scala 29:58]
  wire [7:0] _GEN_824 = 8'ha4 == _T_4[7:0] ? 8'h0 : _GEN_823; // @[Cat.scala 29:58]
  wire [7:0] _GEN_825 = 8'ha5 == _T_4[7:0] ? 8'h0 : _GEN_824; // @[Cat.scala 29:58]
  wire [7:0] _GEN_826 = 8'ha6 == _T_4[7:0] ? 8'h0 : _GEN_825; // @[Cat.scala 29:58]
  wire [7:0] _GEN_827 = 8'ha7 == _T_4[7:0] ? 8'h0 : _GEN_826; // @[Cat.scala 29:58]
  wire [7:0] _GEN_828 = 8'ha8 == _T_4[7:0] ? 8'h0 : _GEN_827; // @[Cat.scala 29:58]
  wire [7:0] _GEN_829 = 8'ha9 == _T_4[7:0] ? 8'h0 : _GEN_828; // @[Cat.scala 29:58]
  wire [7:0] _GEN_830 = 8'haa == _T_4[7:0] ? 8'h0 : _GEN_829; // @[Cat.scala 29:58]
  wire [7:0] _GEN_831 = 8'hab == _T_4[7:0] ? 8'h0 : _GEN_830; // @[Cat.scala 29:58]
  wire [7:0] _GEN_832 = 8'hac == _T_4[7:0] ? 8'h0 : _GEN_831; // @[Cat.scala 29:58]
  wire [7:0] _GEN_833 = 8'had == _T_4[7:0] ? 8'h0 : _GEN_832; // @[Cat.scala 29:58]
  wire [7:0] _GEN_834 = 8'hae == _T_4[7:0] ? 8'h0 : _GEN_833; // @[Cat.scala 29:58]
  wire [7:0] _GEN_835 = 8'haf == _T_4[7:0] ? 8'h0 : _GEN_834; // @[Cat.scala 29:58]
  wire [7:0] _GEN_836 = 8'hb0 == _T_4[7:0] ? 8'h0 : _GEN_835; // @[Cat.scala 29:58]
  wire [7:0] _GEN_837 = 8'hb1 == _T_4[7:0] ? 8'h0 : _GEN_836; // @[Cat.scala 29:58]
  wire [7:0] _GEN_838 = 8'hb2 == _T_4[7:0] ? 8'h0 : _GEN_837; // @[Cat.scala 29:58]
  wire [7:0] _GEN_839 = 8'hb3 == _T_4[7:0] ? 8'h0 : _GEN_838; // @[Cat.scala 29:58]
  wire [7:0] _GEN_840 = 8'hb4 == _T_4[7:0] ? 8'h0 : _GEN_839; // @[Cat.scala 29:58]
  wire [7:0] _GEN_841 = 8'hb5 == _T_4[7:0] ? 8'h0 : _GEN_840; // @[Cat.scala 29:58]
  wire [7:0] _GEN_842 = 8'hb6 == _T_4[7:0] ? 8'h0 : _GEN_841; // @[Cat.scala 29:58]
  wire [7:0] _GEN_843 = 8'hb7 == _T_4[7:0] ? 8'h0 : _GEN_842; // @[Cat.scala 29:58]
  wire [7:0] _GEN_844 = 8'hb8 == _T_4[7:0] ? 8'h0 : _GEN_843; // @[Cat.scala 29:58]
  wire [7:0] _GEN_845 = 8'hb9 == _T_4[7:0] ? 8'h0 : _GEN_844; // @[Cat.scala 29:58]
  wire [7:0] _GEN_846 = 8'hba == _T_4[7:0] ? 8'h0 : _GEN_845; // @[Cat.scala 29:58]
  wire [7:0] _GEN_847 = 8'hbb == _T_4[7:0] ? 8'h0 : _GEN_846; // @[Cat.scala 29:58]
  wire [7:0] _GEN_848 = 8'hbc == _T_4[7:0] ? 8'h0 : _GEN_847; // @[Cat.scala 29:58]
  wire [7:0] _GEN_849 = 8'hbd == _T_4[7:0] ? 8'h0 : _GEN_848; // @[Cat.scala 29:58]
  wire [7:0] _GEN_850 = 8'hbe == _T_4[7:0] ? 8'h0 : _GEN_849; // @[Cat.scala 29:58]
  wire [7:0] _GEN_851 = 8'hbf == _T_4[7:0] ? 8'h0 : _GEN_850; // @[Cat.scala 29:58]
  wire [7:0] _GEN_852 = 8'hc0 == _T_4[7:0] ? 8'h0 : _GEN_851; // @[Cat.scala 29:58]
  wire [7:0] _GEN_853 = 8'hc1 == _T_4[7:0] ? 8'h0 : _GEN_852; // @[Cat.scala 29:58]
  wire [7:0] _GEN_854 = 8'hc2 == _T_4[7:0] ? 8'h0 : _GEN_853; // @[Cat.scala 29:58]
  wire [7:0] _GEN_855 = 8'hc3 == _T_4[7:0] ? 8'h0 : _GEN_854; // @[Cat.scala 29:58]
  wire [7:0] _GEN_856 = 8'hc4 == _T_4[7:0] ? 8'h0 : _GEN_855; // @[Cat.scala 29:58]
  wire [7:0] _GEN_857 = 8'hc5 == _T_4[7:0] ? 8'h0 : _GEN_856; // @[Cat.scala 29:58]
  wire [7:0] _GEN_858 = 8'hc6 == _T_4[7:0] ? 8'h0 : _GEN_857; // @[Cat.scala 29:58]
  wire [7:0] _GEN_859 = 8'hc7 == _T_4[7:0] ? 8'h0 : _GEN_858; // @[Cat.scala 29:58]
  wire [7:0] _GEN_860 = 8'hc8 == _T_4[7:0] ? 8'h0 : _GEN_859; // @[Cat.scala 29:58]
  wire [7:0] _GEN_861 = 8'hc9 == _T_4[7:0] ? 8'h0 : _GEN_860; // @[Cat.scala 29:58]
  wire [7:0] _GEN_862 = 8'hca == _T_4[7:0] ? 8'h0 : _GEN_861; // @[Cat.scala 29:58]
  wire [7:0] _GEN_863 = 8'hcb == _T_4[7:0] ? 8'h0 : _GEN_862; // @[Cat.scala 29:58]
  wire [7:0] _GEN_864 = 8'hcc == _T_4[7:0] ? 8'h0 : _GEN_863; // @[Cat.scala 29:58]
  wire [7:0] _GEN_865 = 8'hcd == _T_4[7:0] ? 8'h0 : _GEN_864; // @[Cat.scala 29:58]
  wire [7:0] _GEN_866 = 8'hce == _T_4[7:0] ? 8'h0 : _GEN_865; // @[Cat.scala 29:58]
  wire [7:0] _GEN_867 = 8'hcf == _T_4[7:0] ? 8'h0 : _GEN_866; // @[Cat.scala 29:58]
  wire [7:0] _GEN_868 = 8'hd0 == _T_4[7:0] ? 8'h0 : _GEN_867; // @[Cat.scala 29:58]
  wire [7:0] _GEN_869 = 8'hd1 == _T_4[7:0] ? 8'h0 : _GEN_868; // @[Cat.scala 29:58]
  wire [7:0] _GEN_870 = 8'hd2 == _T_4[7:0] ? 8'h0 : _GEN_869; // @[Cat.scala 29:58]
  wire [7:0] _GEN_871 = 8'hd3 == _T_4[7:0] ? 8'h0 : _GEN_870; // @[Cat.scala 29:58]
  wire [7:0] _GEN_872 = 8'hd4 == _T_4[7:0] ? 8'h0 : _GEN_871; // @[Cat.scala 29:58]
  wire [7:0] _GEN_873 = 8'hd5 == _T_4[7:0] ? 8'h0 : _GEN_872; // @[Cat.scala 29:58]
  wire [7:0] _GEN_874 = 8'hd6 == _T_4[7:0] ? 8'h0 : _GEN_873; // @[Cat.scala 29:58]
  wire [7:0] _GEN_875 = 8'hd7 == _T_4[7:0] ? 8'h0 : _GEN_874; // @[Cat.scala 29:58]
  wire [7:0] _GEN_876 = 8'hd8 == _T_4[7:0] ? 8'h0 : _GEN_875; // @[Cat.scala 29:58]
  wire [7:0] _GEN_877 = 8'hd9 == _T_4[7:0] ? 8'h0 : _GEN_876; // @[Cat.scala 29:58]
  wire [7:0] _GEN_878 = 8'hda == _T_4[7:0] ? 8'h0 : _GEN_877; // @[Cat.scala 29:58]
  wire [7:0] _GEN_879 = 8'hdb == _T_4[7:0] ? 8'h0 : _GEN_878; // @[Cat.scala 29:58]
  wire [15:0] _T_11 = {_GEN_659,_GEN_879}; // @[Cat.scala 29:58]
  reg [31:0] addr; // @[ROM.scala 26:21]
  reg  _T_14; // @[ROM.scala 28:15]
  wire [31:0] _T_16 = addr + 32'h3; // @[ROM.scala 29:40]
  wire [31:0] _T_20 = addr + 32'h2; // @[ROM.scala 29:58]
  wire [31:0] _T_24 = addr + 32'h1; // @[ROM.scala 29:76]
  wire [7:0] _GEN_881 = 8'h1 == _T_24[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_882 = 8'h2 == _T_24[7:0] ? 8'h0 : _GEN_881; // @[Cat.scala 29:58]
  wire [7:0] _GEN_883 = 8'h3 == _T_24[7:0] ? 8'hfe : _GEN_882; // @[Cat.scala 29:58]
  wire [7:0] _GEN_884 = 8'h4 == _T_24[7:0] ? 8'h93 : _GEN_883; // @[Cat.scala 29:58]
  wire [7:0] _GEN_885 = 8'h5 == _T_24[7:0] ? 8'h5 : _GEN_884; // @[Cat.scala 29:58]
  wire [7:0] _GEN_886 = 8'h6 == _T_24[7:0] ? 8'h0 : _GEN_885; // @[Cat.scala 29:58]
  wire [7:0] _GEN_887 = 8'h7 == _T_24[7:0] ? 8'hfc : _GEN_886; // @[Cat.scala 29:58]
  wire [7:0] _GEN_888 = 8'h8 == _T_24[7:0] ? 8'h33 : _GEN_887; // @[Cat.scala 29:58]
  wire [7:0] _GEN_889 = 8'h9 == _T_24[7:0] ? 8'h6 : _GEN_888; // @[Cat.scala 29:58]
  wire [7:0] _GEN_890 = 8'ha == _T_24[7:0] ? 8'hb5 : _GEN_889; // @[Cat.scala 29:58]
  wire [7:0] _GEN_891 = 8'hb == _T_24[7:0] ? 8'h0 : _GEN_890; // @[Cat.scala 29:58]
  wire [7:0] _GEN_892 = 8'hc == _T_24[7:0] ? 8'h13 : _GEN_891; // @[Cat.scala 29:58]
  wire [7:0] _GEN_893 = 8'hd == _T_24[7:0] ? 8'h5 : _GEN_892; // @[Cat.scala 29:58]
  wire [7:0] _GEN_894 = 8'he == _T_24[7:0] ? 8'ha0 : _GEN_893; // @[Cat.scala 29:58]
  wire [7:0] _GEN_895 = 8'hf == _T_24[7:0] ? 8'h0 : _GEN_894; // @[Cat.scala 29:58]
  wire [7:0] _GEN_896 = 8'h10 == _T_24[7:0] ? 8'h73 : _GEN_895; // @[Cat.scala 29:58]
  wire [7:0] _GEN_897 = 8'h11 == _T_24[7:0] ? 8'h0 : _GEN_896; // @[Cat.scala 29:58]
  wire [7:0] _GEN_898 = 8'h12 == _T_24[7:0] ? 8'h0 : _GEN_897; // @[Cat.scala 29:58]
  wire [7:0] _GEN_899 = 8'h13 == _T_24[7:0] ? 8'h0 : _GEN_898; // @[Cat.scala 29:58]
  wire [7:0] _GEN_900 = 8'h14 == _T_24[7:0] ? 8'h0 : _GEN_899; // @[Cat.scala 29:58]
  wire [7:0] _GEN_901 = 8'h15 == _T_24[7:0] ? 8'h0 : _GEN_900; // @[Cat.scala 29:58]
  wire [7:0] _GEN_902 = 8'h16 == _T_24[7:0] ? 8'h0 : _GEN_901; // @[Cat.scala 29:58]
  wire [7:0] _GEN_903 = 8'h17 == _T_24[7:0] ? 8'h0 : _GEN_902; // @[Cat.scala 29:58]
  wire [7:0] _GEN_904 = 8'h18 == _T_24[7:0] ? 8'h0 : _GEN_903; // @[Cat.scala 29:58]
  wire [7:0] _GEN_905 = 8'h19 == _T_24[7:0] ? 8'h0 : _GEN_904; // @[Cat.scala 29:58]
  wire [7:0] _GEN_906 = 8'h1a == _T_24[7:0] ? 8'h0 : _GEN_905; // @[Cat.scala 29:58]
  wire [7:0] _GEN_907 = 8'h1b == _T_24[7:0] ? 8'h0 : _GEN_906; // @[Cat.scala 29:58]
  wire [7:0] _GEN_908 = 8'h1c == _T_24[7:0] ? 8'h0 : _GEN_907; // @[Cat.scala 29:58]
  wire [7:0] _GEN_909 = 8'h1d == _T_24[7:0] ? 8'h0 : _GEN_908; // @[Cat.scala 29:58]
  wire [7:0] _GEN_910 = 8'h1e == _T_24[7:0] ? 8'h0 : _GEN_909; // @[Cat.scala 29:58]
  wire [7:0] _GEN_911 = 8'h1f == _T_24[7:0] ? 8'h0 : _GEN_910; // @[Cat.scala 29:58]
  wire [7:0] _GEN_912 = 8'h20 == _T_24[7:0] ? 8'h0 : _GEN_911; // @[Cat.scala 29:58]
  wire [7:0] _GEN_913 = 8'h21 == _T_24[7:0] ? 8'h0 : _GEN_912; // @[Cat.scala 29:58]
  wire [7:0] _GEN_914 = 8'h22 == _T_24[7:0] ? 8'h0 : _GEN_913; // @[Cat.scala 29:58]
  wire [7:0] _GEN_915 = 8'h23 == _T_24[7:0] ? 8'h0 : _GEN_914; // @[Cat.scala 29:58]
  wire [7:0] _GEN_916 = 8'h24 == _T_24[7:0] ? 8'h0 : _GEN_915; // @[Cat.scala 29:58]
  wire [7:0] _GEN_917 = 8'h25 == _T_24[7:0] ? 8'h0 : _GEN_916; // @[Cat.scala 29:58]
  wire [7:0] _GEN_918 = 8'h26 == _T_24[7:0] ? 8'h0 : _GEN_917; // @[Cat.scala 29:58]
  wire [7:0] _GEN_919 = 8'h27 == _T_24[7:0] ? 8'h0 : _GEN_918; // @[Cat.scala 29:58]
  wire [7:0] _GEN_920 = 8'h28 == _T_24[7:0] ? 8'h0 : _GEN_919; // @[Cat.scala 29:58]
  wire [7:0] _GEN_921 = 8'h29 == _T_24[7:0] ? 8'h0 : _GEN_920; // @[Cat.scala 29:58]
  wire [7:0] _GEN_922 = 8'h2a == _T_24[7:0] ? 8'h0 : _GEN_921; // @[Cat.scala 29:58]
  wire [7:0] _GEN_923 = 8'h2b == _T_24[7:0] ? 8'h0 : _GEN_922; // @[Cat.scala 29:58]
  wire [7:0] _GEN_924 = 8'h2c == _T_24[7:0] ? 8'h0 : _GEN_923; // @[Cat.scala 29:58]
  wire [7:0] _GEN_925 = 8'h2d == _T_24[7:0] ? 8'h0 : _GEN_924; // @[Cat.scala 29:58]
  wire [7:0] _GEN_926 = 8'h2e == _T_24[7:0] ? 8'h0 : _GEN_925; // @[Cat.scala 29:58]
  wire [7:0] _GEN_927 = 8'h2f == _T_24[7:0] ? 8'h0 : _GEN_926; // @[Cat.scala 29:58]
  wire [7:0] _GEN_928 = 8'h30 == _T_24[7:0] ? 8'h0 : _GEN_927; // @[Cat.scala 29:58]
  wire [7:0] _GEN_929 = 8'h31 == _T_24[7:0] ? 8'h0 : _GEN_928; // @[Cat.scala 29:58]
  wire [7:0] _GEN_930 = 8'h32 == _T_24[7:0] ? 8'h0 : _GEN_929; // @[Cat.scala 29:58]
  wire [7:0] _GEN_931 = 8'h33 == _T_24[7:0] ? 8'h0 : _GEN_930; // @[Cat.scala 29:58]
  wire [7:0] _GEN_932 = 8'h34 == _T_24[7:0] ? 8'h0 : _GEN_931; // @[Cat.scala 29:58]
  wire [7:0] _GEN_933 = 8'h35 == _T_24[7:0] ? 8'h0 : _GEN_932; // @[Cat.scala 29:58]
  wire [7:0] _GEN_934 = 8'h36 == _T_24[7:0] ? 8'h0 : _GEN_933; // @[Cat.scala 29:58]
  wire [7:0] _GEN_935 = 8'h37 == _T_24[7:0] ? 8'h0 : _GEN_934; // @[Cat.scala 29:58]
  wire [7:0] _GEN_936 = 8'h38 == _T_24[7:0] ? 8'h0 : _GEN_935; // @[Cat.scala 29:58]
  wire [7:0] _GEN_937 = 8'h39 == _T_24[7:0] ? 8'h0 : _GEN_936; // @[Cat.scala 29:58]
  wire [7:0] _GEN_938 = 8'h3a == _T_24[7:0] ? 8'h0 : _GEN_937; // @[Cat.scala 29:58]
  wire [7:0] _GEN_939 = 8'h3b == _T_24[7:0] ? 8'h0 : _GEN_938; // @[Cat.scala 29:58]
  wire [7:0] _GEN_940 = 8'h3c == _T_24[7:0] ? 8'h0 : _GEN_939; // @[Cat.scala 29:58]
  wire [7:0] _GEN_941 = 8'h3d == _T_24[7:0] ? 8'h0 : _GEN_940; // @[Cat.scala 29:58]
  wire [7:0] _GEN_942 = 8'h3e == _T_24[7:0] ? 8'h0 : _GEN_941; // @[Cat.scala 29:58]
  wire [7:0] _GEN_943 = 8'h3f == _T_24[7:0] ? 8'h0 : _GEN_942; // @[Cat.scala 29:58]
  wire [7:0] _GEN_944 = 8'h40 == _T_24[7:0] ? 8'h0 : _GEN_943; // @[Cat.scala 29:58]
  wire [7:0] _GEN_945 = 8'h41 == _T_24[7:0] ? 8'h0 : _GEN_944; // @[Cat.scala 29:58]
  wire [7:0] _GEN_946 = 8'h42 == _T_24[7:0] ? 8'h0 : _GEN_945; // @[Cat.scala 29:58]
  wire [7:0] _GEN_947 = 8'h43 == _T_24[7:0] ? 8'h0 : _GEN_946; // @[Cat.scala 29:58]
  wire [7:0] _GEN_948 = 8'h44 == _T_24[7:0] ? 8'h0 : _GEN_947; // @[Cat.scala 29:58]
  wire [7:0] _GEN_949 = 8'h45 == _T_24[7:0] ? 8'h0 : _GEN_948; // @[Cat.scala 29:58]
  wire [7:0] _GEN_950 = 8'h46 == _T_24[7:0] ? 8'h0 : _GEN_949; // @[Cat.scala 29:58]
  wire [7:0] _GEN_951 = 8'h47 == _T_24[7:0] ? 8'h0 : _GEN_950; // @[Cat.scala 29:58]
  wire [7:0] _GEN_952 = 8'h48 == _T_24[7:0] ? 8'h0 : _GEN_951; // @[Cat.scala 29:58]
  wire [7:0] _GEN_953 = 8'h49 == _T_24[7:0] ? 8'h0 : _GEN_952; // @[Cat.scala 29:58]
  wire [7:0] _GEN_954 = 8'h4a == _T_24[7:0] ? 8'h0 : _GEN_953; // @[Cat.scala 29:58]
  wire [7:0] _GEN_955 = 8'h4b == _T_24[7:0] ? 8'h0 : _GEN_954; // @[Cat.scala 29:58]
  wire [7:0] _GEN_956 = 8'h4c == _T_24[7:0] ? 8'h0 : _GEN_955; // @[Cat.scala 29:58]
  wire [7:0] _GEN_957 = 8'h4d == _T_24[7:0] ? 8'h0 : _GEN_956; // @[Cat.scala 29:58]
  wire [7:0] _GEN_958 = 8'h4e == _T_24[7:0] ? 8'h0 : _GEN_957; // @[Cat.scala 29:58]
  wire [7:0] _GEN_959 = 8'h4f == _T_24[7:0] ? 8'h0 : _GEN_958; // @[Cat.scala 29:58]
  wire [7:0] _GEN_960 = 8'h50 == _T_24[7:0] ? 8'h0 : _GEN_959; // @[Cat.scala 29:58]
  wire [7:0] _GEN_961 = 8'h51 == _T_24[7:0] ? 8'h0 : _GEN_960; // @[Cat.scala 29:58]
  wire [7:0] _GEN_962 = 8'h52 == _T_24[7:0] ? 8'h0 : _GEN_961; // @[Cat.scala 29:58]
  wire [7:0] _GEN_963 = 8'h53 == _T_24[7:0] ? 8'h0 : _GEN_962; // @[Cat.scala 29:58]
  wire [7:0] _GEN_964 = 8'h54 == _T_24[7:0] ? 8'h0 : _GEN_963; // @[Cat.scala 29:58]
  wire [7:0] _GEN_965 = 8'h55 == _T_24[7:0] ? 8'h0 : _GEN_964; // @[Cat.scala 29:58]
  wire [7:0] _GEN_966 = 8'h56 == _T_24[7:0] ? 8'h0 : _GEN_965; // @[Cat.scala 29:58]
  wire [7:0] _GEN_967 = 8'h57 == _T_24[7:0] ? 8'h0 : _GEN_966; // @[Cat.scala 29:58]
  wire [7:0] _GEN_968 = 8'h58 == _T_24[7:0] ? 8'h0 : _GEN_967; // @[Cat.scala 29:58]
  wire [7:0] _GEN_969 = 8'h59 == _T_24[7:0] ? 8'h0 : _GEN_968; // @[Cat.scala 29:58]
  wire [7:0] _GEN_970 = 8'h5a == _T_24[7:0] ? 8'h0 : _GEN_969; // @[Cat.scala 29:58]
  wire [7:0] _GEN_971 = 8'h5b == _T_24[7:0] ? 8'h0 : _GEN_970; // @[Cat.scala 29:58]
  wire [7:0] _GEN_972 = 8'h5c == _T_24[7:0] ? 8'h0 : _GEN_971; // @[Cat.scala 29:58]
  wire [7:0] _GEN_973 = 8'h5d == _T_24[7:0] ? 8'h0 : _GEN_972; // @[Cat.scala 29:58]
  wire [7:0] _GEN_974 = 8'h5e == _T_24[7:0] ? 8'h0 : _GEN_973; // @[Cat.scala 29:58]
  wire [7:0] _GEN_975 = 8'h5f == _T_24[7:0] ? 8'h0 : _GEN_974; // @[Cat.scala 29:58]
  wire [7:0] _GEN_976 = 8'h60 == _T_24[7:0] ? 8'h0 : _GEN_975; // @[Cat.scala 29:58]
  wire [7:0] _GEN_977 = 8'h61 == _T_24[7:0] ? 8'h0 : _GEN_976; // @[Cat.scala 29:58]
  wire [7:0] _GEN_978 = 8'h62 == _T_24[7:0] ? 8'h0 : _GEN_977; // @[Cat.scala 29:58]
  wire [7:0] _GEN_979 = 8'h63 == _T_24[7:0] ? 8'h0 : _GEN_978; // @[Cat.scala 29:58]
  wire [7:0] _GEN_980 = 8'h64 == _T_24[7:0] ? 8'h0 : _GEN_979; // @[Cat.scala 29:58]
  wire [7:0] _GEN_981 = 8'h65 == _T_24[7:0] ? 8'h0 : _GEN_980; // @[Cat.scala 29:58]
  wire [7:0] _GEN_982 = 8'h66 == _T_24[7:0] ? 8'h0 : _GEN_981; // @[Cat.scala 29:58]
  wire [7:0] _GEN_983 = 8'h67 == _T_24[7:0] ? 8'h0 : _GEN_982; // @[Cat.scala 29:58]
  wire [7:0] _GEN_984 = 8'h68 == _T_24[7:0] ? 8'h0 : _GEN_983; // @[Cat.scala 29:58]
  wire [7:0] _GEN_985 = 8'h69 == _T_24[7:0] ? 8'h0 : _GEN_984; // @[Cat.scala 29:58]
  wire [7:0] _GEN_986 = 8'h6a == _T_24[7:0] ? 8'h0 : _GEN_985; // @[Cat.scala 29:58]
  wire [7:0] _GEN_987 = 8'h6b == _T_24[7:0] ? 8'h0 : _GEN_986; // @[Cat.scala 29:58]
  wire [7:0] _GEN_988 = 8'h6c == _T_24[7:0] ? 8'h0 : _GEN_987; // @[Cat.scala 29:58]
  wire [7:0] _GEN_989 = 8'h6d == _T_24[7:0] ? 8'h0 : _GEN_988; // @[Cat.scala 29:58]
  wire [7:0] _GEN_990 = 8'h6e == _T_24[7:0] ? 8'h0 : _GEN_989; // @[Cat.scala 29:58]
  wire [7:0] _GEN_991 = 8'h6f == _T_24[7:0] ? 8'h0 : _GEN_990; // @[Cat.scala 29:58]
  wire [7:0] _GEN_992 = 8'h70 == _T_24[7:0] ? 8'h0 : _GEN_991; // @[Cat.scala 29:58]
  wire [7:0] _GEN_993 = 8'h71 == _T_24[7:0] ? 8'h0 : _GEN_992; // @[Cat.scala 29:58]
  wire [7:0] _GEN_994 = 8'h72 == _T_24[7:0] ? 8'h0 : _GEN_993; // @[Cat.scala 29:58]
  wire [7:0] _GEN_995 = 8'h73 == _T_24[7:0] ? 8'h0 : _GEN_994; // @[Cat.scala 29:58]
  wire [7:0] _GEN_996 = 8'h74 == _T_24[7:0] ? 8'h0 : _GEN_995; // @[Cat.scala 29:58]
  wire [7:0] _GEN_997 = 8'h75 == _T_24[7:0] ? 8'h0 : _GEN_996; // @[Cat.scala 29:58]
  wire [7:0] _GEN_998 = 8'h76 == _T_24[7:0] ? 8'h0 : _GEN_997; // @[Cat.scala 29:58]
  wire [7:0] _GEN_999 = 8'h77 == _T_24[7:0] ? 8'h0 : _GEN_998; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1000 = 8'h78 == _T_24[7:0] ? 8'h0 : _GEN_999; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1001 = 8'h79 == _T_24[7:0] ? 8'h0 : _GEN_1000; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1002 = 8'h7a == _T_24[7:0] ? 8'h0 : _GEN_1001; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1003 = 8'h7b == _T_24[7:0] ? 8'h0 : _GEN_1002; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1004 = 8'h7c == _T_24[7:0] ? 8'h0 : _GEN_1003; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1005 = 8'h7d == _T_24[7:0] ? 8'h0 : _GEN_1004; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1006 = 8'h7e == _T_24[7:0] ? 8'h0 : _GEN_1005; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1007 = 8'h7f == _T_24[7:0] ? 8'h0 : _GEN_1006; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1008 = 8'h80 == _T_24[7:0] ? 8'h0 : _GEN_1007; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1009 = 8'h81 == _T_24[7:0] ? 8'h0 : _GEN_1008; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1010 = 8'h82 == _T_24[7:0] ? 8'h0 : _GEN_1009; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1011 = 8'h83 == _T_24[7:0] ? 8'h0 : _GEN_1010; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1012 = 8'h84 == _T_24[7:0] ? 8'h0 : _GEN_1011; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1013 = 8'h85 == _T_24[7:0] ? 8'h0 : _GEN_1012; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1014 = 8'h86 == _T_24[7:0] ? 8'h0 : _GEN_1013; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1015 = 8'h87 == _T_24[7:0] ? 8'h0 : _GEN_1014; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1016 = 8'h88 == _T_24[7:0] ? 8'h0 : _GEN_1015; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1017 = 8'h89 == _T_24[7:0] ? 8'h0 : _GEN_1016; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1018 = 8'h8a == _T_24[7:0] ? 8'h0 : _GEN_1017; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1019 = 8'h8b == _T_24[7:0] ? 8'h0 : _GEN_1018; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1020 = 8'h8c == _T_24[7:0] ? 8'h0 : _GEN_1019; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1021 = 8'h8d == _T_24[7:0] ? 8'h0 : _GEN_1020; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1022 = 8'h8e == _T_24[7:0] ? 8'h0 : _GEN_1021; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1023 = 8'h8f == _T_24[7:0] ? 8'h0 : _GEN_1022; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1024 = 8'h90 == _T_24[7:0] ? 8'h0 : _GEN_1023; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1025 = 8'h91 == _T_24[7:0] ? 8'h0 : _GEN_1024; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1026 = 8'h92 == _T_24[7:0] ? 8'h0 : _GEN_1025; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1027 = 8'h93 == _T_24[7:0] ? 8'h0 : _GEN_1026; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1028 = 8'h94 == _T_24[7:0] ? 8'h0 : _GEN_1027; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1029 = 8'h95 == _T_24[7:0] ? 8'h0 : _GEN_1028; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1030 = 8'h96 == _T_24[7:0] ? 8'h0 : _GEN_1029; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1031 = 8'h97 == _T_24[7:0] ? 8'h0 : _GEN_1030; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1032 = 8'h98 == _T_24[7:0] ? 8'h0 : _GEN_1031; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1033 = 8'h99 == _T_24[7:0] ? 8'h0 : _GEN_1032; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1034 = 8'h9a == _T_24[7:0] ? 8'h0 : _GEN_1033; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1035 = 8'h9b == _T_24[7:0] ? 8'h0 : _GEN_1034; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1036 = 8'h9c == _T_24[7:0] ? 8'h0 : _GEN_1035; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1037 = 8'h9d == _T_24[7:0] ? 8'h0 : _GEN_1036; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1038 = 8'h9e == _T_24[7:0] ? 8'h0 : _GEN_1037; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1039 = 8'h9f == _T_24[7:0] ? 8'h0 : _GEN_1038; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1040 = 8'ha0 == _T_24[7:0] ? 8'h0 : _GEN_1039; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1041 = 8'ha1 == _T_24[7:0] ? 8'h0 : _GEN_1040; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1042 = 8'ha2 == _T_24[7:0] ? 8'h0 : _GEN_1041; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1043 = 8'ha3 == _T_24[7:0] ? 8'h0 : _GEN_1042; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1044 = 8'ha4 == _T_24[7:0] ? 8'h0 : _GEN_1043; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1045 = 8'ha5 == _T_24[7:0] ? 8'h0 : _GEN_1044; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1046 = 8'ha6 == _T_24[7:0] ? 8'h0 : _GEN_1045; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1047 = 8'ha7 == _T_24[7:0] ? 8'h0 : _GEN_1046; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1048 = 8'ha8 == _T_24[7:0] ? 8'h0 : _GEN_1047; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1049 = 8'ha9 == _T_24[7:0] ? 8'h0 : _GEN_1048; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1050 = 8'haa == _T_24[7:0] ? 8'h0 : _GEN_1049; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1051 = 8'hab == _T_24[7:0] ? 8'h0 : _GEN_1050; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1052 = 8'hac == _T_24[7:0] ? 8'h0 : _GEN_1051; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1053 = 8'had == _T_24[7:0] ? 8'h0 : _GEN_1052; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1054 = 8'hae == _T_24[7:0] ? 8'h0 : _GEN_1053; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1055 = 8'haf == _T_24[7:0] ? 8'h0 : _GEN_1054; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1056 = 8'hb0 == _T_24[7:0] ? 8'h0 : _GEN_1055; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1057 = 8'hb1 == _T_24[7:0] ? 8'h0 : _GEN_1056; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1058 = 8'hb2 == _T_24[7:0] ? 8'h0 : _GEN_1057; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1059 = 8'hb3 == _T_24[7:0] ? 8'h0 : _GEN_1058; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1060 = 8'hb4 == _T_24[7:0] ? 8'h0 : _GEN_1059; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1061 = 8'hb5 == _T_24[7:0] ? 8'h0 : _GEN_1060; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1062 = 8'hb6 == _T_24[7:0] ? 8'h0 : _GEN_1061; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1063 = 8'hb7 == _T_24[7:0] ? 8'h0 : _GEN_1062; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1064 = 8'hb8 == _T_24[7:0] ? 8'h0 : _GEN_1063; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1065 = 8'hb9 == _T_24[7:0] ? 8'h0 : _GEN_1064; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1066 = 8'hba == _T_24[7:0] ? 8'h0 : _GEN_1065; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1067 = 8'hbb == _T_24[7:0] ? 8'h0 : _GEN_1066; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1068 = 8'hbc == _T_24[7:0] ? 8'h0 : _GEN_1067; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1069 = 8'hbd == _T_24[7:0] ? 8'h0 : _GEN_1068; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1070 = 8'hbe == _T_24[7:0] ? 8'h0 : _GEN_1069; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1071 = 8'hbf == _T_24[7:0] ? 8'h0 : _GEN_1070; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1072 = 8'hc0 == _T_24[7:0] ? 8'h0 : _GEN_1071; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1073 = 8'hc1 == _T_24[7:0] ? 8'h0 : _GEN_1072; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1074 = 8'hc2 == _T_24[7:0] ? 8'h0 : _GEN_1073; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1075 = 8'hc3 == _T_24[7:0] ? 8'h0 : _GEN_1074; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1076 = 8'hc4 == _T_24[7:0] ? 8'h0 : _GEN_1075; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1077 = 8'hc5 == _T_24[7:0] ? 8'h0 : _GEN_1076; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1078 = 8'hc6 == _T_24[7:0] ? 8'h0 : _GEN_1077; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1079 = 8'hc7 == _T_24[7:0] ? 8'h0 : _GEN_1078; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1080 = 8'hc8 == _T_24[7:0] ? 8'h0 : _GEN_1079; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1081 = 8'hc9 == _T_24[7:0] ? 8'h0 : _GEN_1080; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1082 = 8'hca == _T_24[7:0] ? 8'h0 : _GEN_1081; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1083 = 8'hcb == _T_24[7:0] ? 8'h0 : _GEN_1082; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1084 = 8'hcc == _T_24[7:0] ? 8'h0 : _GEN_1083; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1085 = 8'hcd == _T_24[7:0] ? 8'h0 : _GEN_1084; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1086 = 8'hce == _T_24[7:0] ? 8'h0 : _GEN_1085; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1087 = 8'hcf == _T_24[7:0] ? 8'h0 : _GEN_1086; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1088 = 8'hd0 == _T_24[7:0] ? 8'h0 : _GEN_1087; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1089 = 8'hd1 == _T_24[7:0] ? 8'h0 : _GEN_1088; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1090 = 8'hd2 == _T_24[7:0] ? 8'h0 : _GEN_1089; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1091 = 8'hd3 == _T_24[7:0] ? 8'h0 : _GEN_1090; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1092 = 8'hd4 == _T_24[7:0] ? 8'h0 : _GEN_1091; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1093 = 8'hd5 == _T_24[7:0] ? 8'h0 : _GEN_1092; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1094 = 8'hd6 == _T_24[7:0] ? 8'h0 : _GEN_1093; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1095 = 8'hd7 == _T_24[7:0] ? 8'h0 : _GEN_1094; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1096 = 8'hd8 == _T_24[7:0] ? 8'h0 : _GEN_1095; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1097 = 8'hd9 == _T_24[7:0] ? 8'h0 : _GEN_1096; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1098 = 8'hda == _T_24[7:0] ? 8'h0 : _GEN_1097; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1099 = 8'hdb == _T_24[7:0] ? 8'h0 : _GEN_1098; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1101 = 8'h1 == addr[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1102 = 8'h2 == addr[7:0] ? 8'h0 : _GEN_1101; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1103 = 8'h3 == addr[7:0] ? 8'hfe : _GEN_1102; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1104 = 8'h4 == addr[7:0] ? 8'h93 : _GEN_1103; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1105 = 8'h5 == addr[7:0] ? 8'h5 : _GEN_1104; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1106 = 8'h6 == addr[7:0] ? 8'h0 : _GEN_1105; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1107 = 8'h7 == addr[7:0] ? 8'hfc : _GEN_1106; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1108 = 8'h8 == addr[7:0] ? 8'h33 : _GEN_1107; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1109 = 8'h9 == addr[7:0] ? 8'h6 : _GEN_1108; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1110 = 8'ha == addr[7:0] ? 8'hb5 : _GEN_1109; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1111 = 8'hb == addr[7:0] ? 8'h0 : _GEN_1110; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1112 = 8'hc == addr[7:0] ? 8'h13 : _GEN_1111; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1113 = 8'hd == addr[7:0] ? 8'h5 : _GEN_1112; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1114 = 8'he == addr[7:0] ? 8'ha0 : _GEN_1113; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1115 = 8'hf == addr[7:0] ? 8'h0 : _GEN_1114; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1116 = 8'h10 == addr[7:0] ? 8'h73 : _GEN_1115; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1117 = 8'h11 == addr[7:0] ? 8'h0 : _GEN_1116; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1118 = 8'h12 == addr[7:0] ? 8'h0 : _GEN_1117; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1119 = 8'h13 == addr[7:0] ? 8'h0 : _GEN_1118; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1120 = 8'h14 == addr[7:0] ? 8'h0 : _GEN_1119; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1121 = 8'h15 == addr[7:0] ? 8'h0 : _GEN_1120; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1122 = 8'h16 == addr[7:0] ? 8'h0 : _GEN_1121; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1123 = 8'h17 == addr[7:0] ? 8'h0 : _GEN_1122; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1124 = 8'h18 == addr[7:0] ? 8'h0 : _GEN_1123; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1125 = 8'h19 == addr[7:0] ? 8'h0 : _GEN_1124; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1126 = 8'h1a == addr[7:0] ? 8'h0 : _GEN_1125; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1127 = 8'h1b == addr[7:0] ? 8'h0 : _GEN_1126; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1128 = 8'h1c == addr[7:0] ? 8'h0 : _GEN_1127; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1129 = 8'h1d == addr[7:0] ? 8'h0 : _GEN_1128; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1130 = 8'h1e == addr[7:0] ? 8'h0 : _GEN_1129; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1131 = 8'h1f == addr[7:0] ? 8'h0 : _GEN_1130; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1132 = 8'h20 == addr[7:0] ? 8'h0 : _GEN_1131; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1133 = 8'h21 == addr[7:0] ? 8'h0 : _GEN_1132; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1134 = 8'h22 == addr[7:0] ? 8'h0 : _GEN_1133; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1135 = 8'h23 == addr[7:0] ? 8'h0 : _GEN_1134; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1136 = 8'h24 == addr[7:0] ? 8'h0 : _GEN_1135; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1137 = 8'h25 == addr[7:0] ? 8'h0 : _GEN_1136; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1138 = 8'h26 == addr[7:0] ? 8'h0 : _GEN_1137; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1139 = 8'h27 == addr[7:0] ? 8'h0 : _GEN_1138; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1140 = 8'h28 == addr[7:0] ? 8'h0 : _GEN_1139; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1141 = 8'h29 == addr[7:0] ? 8'h0 : _GEN_1140; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1142 = 8'h2a == addr[7:0] ? 8'h0 : _GEN_1141; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1143 = 8'h2b == addr[7:0] ? 8'h0 : _GEN_1142; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1144 = 8'h2c == addr[7:0] ? 8'h0 : _GEN_1143; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1145 = 8'h2d == addr[7:0] ? 8'h0 : _GEN_1144; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1146 = 8'h2e == addr[7:0] ? 8'h0 : _GEN_1145; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1147 = 8'h2f == addr[7:0] ? 8'h0 : _GEN_1146; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1148 = 8'h30 == addr[7:0] ? 8'h0 : _GEN_1147; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1149 = 8'h31 == addr[7:0] ? 8'h0 : _GEN_1148; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1150 = 8'h32 == addr[7:0] ? 8'h0 : _GEN_1149; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1151 = 8'h33 == addr[7:0] ? 8'h0 : _GEN_1150; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1152 = 8'h34 == addr[7:0] ? 8'h0 : _GEN_1151; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1153 = 8'h35 == addr[7:0] ? 8'h0 : _GEN_1152; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1154 = 8'h36 == addr[7:0] ? 8'h0 : _GEN_1153; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1155 = 8'h37 == addr[7:0] ? 8'h0 : _GEN_1154; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1156 = 8'h38 == addr[7:0] ? 8'h0 : _GEN_1155; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1157 = 8'h39 == addr[7:0] ? 8'h0 : _GEN_1156; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1158 = 8'h3a == addr[7:0] ? 8'h0 : _GEN_1157; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1159 = 8'h3b == addr[7:0] ? 8'h0 : _GEN_1158; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1160 = 8'h3c == addr[7:0] ? 8'h0 : _GEN_1159; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1161 = 8'h3d == addr[7:0] ? 8'h0 : _GEN_1160; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1162 = 8'h3e == addr[7:0] ? 8'h0 : _GEN_1161; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1163 = 8'h3f == addr[7:0] ? 8'h0 : _GEN_1162; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1164 = 8'h40 == addr[7:0] ? 8'h0 : _GEN_1163; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1165 = 8'h41 == addr[7:0] ? 8'h0 : _GEN_1164; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1166 = 8'h42 == addr[7:0] ? 8'h0 : _GEN_1165; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1167 = 8'h43 == addr[7:0] ? 8'h0 : _GEN_1166; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1168 = 8'h44 == addr[7:0] ? 8'h0 : _GEN_1167; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1169 = 8'h45 == addr[7:0] ? 8'h0 : _GEN_1168; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1170 = 8'h46 == addr[7:0] ? 8'h0 : _GEN_1169; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1171 = 8'h47 == addr[7:0] ? 8'h0 : _GEN_1170; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1172 = 8'h48 == addr[7:0] ? 8'h0 : _GEN_1171; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1173 = 8'h49 == addr[7:0] ? 8'h0 : _GEN_1172; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1174 = 8'h4a == addr[7:0] ? 8'h0 : _GEN_1173; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1175 = 8'h4b == addr[7:0] ? 8'h0 : _GEN_1174; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1176 = 8'h4c == addr[7:0] ? 8'h0 : _GEN_1175; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1177 = 8'h4d == addr[7:0] ? 8'h0 : _GEN_1176; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1178 = 8'h4e == addr[7:0] ? 8'h0 : _GEN_1177; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1179 = 8'h4f == addr[7:0] ? 8'h0 : _GEN_1178; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1180 = 8'h50 == addr[7:0] ? 8'h0 : _GEN_1179; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1181 = 8'h51 == addr[7:0] ? 8'h0 : _GEN_1180; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1182 = 8'h52 == addr[7:0] ? 8'h0 : _GEN_1181; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1183 = 8'h53 == addr[7:0] ? 8'h0 : _GEN_1182; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1184 = 8'h54 == addr[7:0] ? 8'h0 : _GEN_1183; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1185 = 8'h55 == addr[7:0] ? 8'h0 : _GEN_1184; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1186 = 8'h56 == addr[7:0] ? 8'h0 : _GEN_1185; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1187 = 8'h57 == addr[7:0] ? 8'h0 : _GEN_1186; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1188 = 8'h58 == addr[7:0] ? 8'h0 : _GEN_1187; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1189 = 8'h59 == addr[7:0] ? 8'h0 : _GEN_1188; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1190 = 8'h5a == addr[7:0] ? 8'h0 : _GEN_1189; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1191 = 8'h5b == addr[7:0] ? 8'h0 : _GEN_1190; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1192 = 8'h5c == addr[7:0] ? 8'h0 : _GEN_1191; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1193 = 8'h5d == addr[7:0] ? 8'h0 : _GEN_1192; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1194 = 8'h5e == addr[7:0] ? 8'h0 : _GEN_1193; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1195 = 8'h5f == addr[7:0] ? 8'h0 : _GEN_1194; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1196 = 8'h60 == addr[7:0] ? 8'h0 : _GEN_1195; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1197 = 8'h61 == addr[7:0] ? 8'h0 : _GEN_1196; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1198 = 8'h62 == addr[7:0] ? 8'h0 : _GEN_1197; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1199 = 8'h63 == addr[7:0] ? 8'h0 : _GEN_1198; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1200 = 8'h64 == addr[7:0] ? 8'h0 : _GEN_1199; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1201 = 8'h65 == addr[7:0] ? 8'h0 : _GEN_1200; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1202 = 8'h66 == addr[7:0] ? 8'h0 : _GEN_1201; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1203 = 8'h67 == addr[7:0] ? 8'h0 : _GEN_1202; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1204 = 8'h68 == addr[7:0] ? 8'h0 : _GEN_1203; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1205 = 8'h69 == addr[7:0] ? 8'h0 : _GEN_1204; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1206 = 8'h6a == addr[7:0] ? 8'h0 : _GEN_1205; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1207 = 8'h6b == addr[7:0] ? 8'h0 : _GEN_1206; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1208 = 8'h6c == addr[7:0] ? 8'h0 : _GEN_1207; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1209 = 8'h6d == addr[7:0] ? 8'h0 : _GEN_1208; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1210 = 8'h6e == addr[7:0] ? 8'h0 : _GEN_1209; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1211 = 8'h6f == addr[7:0] ? 8'h0 : _GEN_1210; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1212 = 8'h70 == addr[7:0] ? 8'h0 : _GEN_1211; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1213 = 8'h71 == addr[7:0] ? 8'h0 : _GEN_1212; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1214 = 8'h72 == addr[7:0] ? 8'h0 : _GEN_1213; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1215 = 8'h73 == addr[7:0] ? 8'h0 : _GEN_1214; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1216 = 8'h74 == addr[7:0] ? 8'h0 : _GEN_1215; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1217 = 8'h75 == addr[7:0] ? 8'h0 : _GEN_1216; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1218 = 8'h76 == addr[7:0] ? 8'h0 : _GEN_1217; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1219 = 8'h77 == addr[7:0] ? 8'h0 : _GEN_1218; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1220 = 8'h78 == addr[7:0] ? 8'h0 : _GEN_1219; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1221 = 8'h79 == addr[7:0] ? 8'h0 : _GEN_1220; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1222 = 8'h7a == addr[7:0] ? 8'h0 : _GEN_1221; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1223 = 8'h7b == addr[7:0] ? 8'h0 : _GEN_1222; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1224 = 8'h7c == addr[7:0] ? 8'h0 : _GEN_1223; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1225 = 8'h7d == addr[7:0] ? 8'h0 : _GEN_1224; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1226 = 8'h7e == addr[7:0] ? 8'h0 : _GEN_1225; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1227 = 8'h7f == addr[7:0] ? 8'h0 : _GEN_1226; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1228 = 8'h80 == addr[7:0] ? 8'h0 : _GEN_1227; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1229 = 8'h81 == addr[7:0] ? 8'h0 : _GEN_1228; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1230 = 8'h82 == addr[7:0] ? 8'h0 : _GEN_1229; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1231 = 8'h83 == addr[7:0] ? 8'h0 : _GEN_1230; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1232 = 8'h84 == addr[7:0] ? 8'h0 : _GEN_1231; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1233 = 8'h85 == addr[7:0] ? 8'h0 : _GEN_1232; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1234 = 8'h86 == addr[7:0] ? 8'h0 : _GEN_1233; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1235 = 8'h87 == addr[7:0] ? 8'h0 : _GEN_1234; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1236 = 8'h88 == addr[7:0] ? 8'h0 : _GEN_1235; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1237 = 8'h89 == addr[7:0] ? 8'h0 : _GEN_1236; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1238 = 8'h8a == addr[7:0] ? 8'h0 : _GEN_1237; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1239 = 8'h8b == addr[7:0] ? 8'h0 : _GEN_1238; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1240 = 8'h8c == addr[7:0] ? 8'h0 : _GEN_1239; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1241 = 8'h8d == addr[7:0] ? 8'h0 : _GEN_1240; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1242 = 8'h8e == addr[7:0] ? 8'h0 : _GEN_1241; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1243 = 8'h8f == addr[7:0] ? 8'h0 : _GEN_1242; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1244 = 8'h90 == addr[7:0] ? 8'h0 : _GEN_1243; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1245 = 8'h91 == addr[7:0] ? 8'h0 : _GEN_1244; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1246 = 8'h92 == addr[7:0] ? 8'h0 : _GEN_1245; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1247 = 8'h93 == addr[7:0] ? 8'h0 : _GEN_1246; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1248 = 8'h94 == addr[7:0] ? 8'h0 : _GEN_1247; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1249 = 8'h95 == addr[7:0] ? 8'h0 : _GEN_1248; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1250 = 8'h96 == addr[7:0] ? 8'h0 : _GEN_1249; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1251 = 8'h97 == addr[7:0] ? 8'h0 : _GEN_1250; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1252 = 8'h98 == addr[7:0] ? 8'h0 : _GEN_1251; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1253 = 8'h99 == addr[7:0] ? 8'h0 : _GEN_1252; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1254 = 8'h9a == addr[7:0] ? 8'h0 : _GEN_1253; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1255 = 8'h9b == addr[7:0] ? 8'h0 : _GEN_1254; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1256 = 8'h9c == addr[7:0] ? 8'h0 : _GEN_1255; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1257 = 8'h9d == addr[7:0] ? 8'h0 : _GEN_1256; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1258 = 8'h9e == addr[7:0] ? 8'h0 : _GEN_1257; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1259 = 8'h9f == addr[7:0] ? 8'h0 : _GEN_1258; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1260 = 8'ha0 == addr[7:0] ? 8'h0 : _GEN_1259; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1261 = 8'ha1 == addr[7:0] ? 8'h0 : _GEN_1260; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1262 = 8'ha2 == addr[7:0] ? 8'h0 : _GEN_1261; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1263 = 8'ha3 == addr[7:0] ? 8'h0 : _GEN_1262; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1264 = 8'ha4 == addr[7:0] ? 8'h0 : _GEN_1263; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1265 = 8'ha5 == addr[7:0] ? 8'h0 : _GEN_1264; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1266 = 8'ha6 == addr[7:0] ? 8'h0 : _GEN_1265; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1267 = 8'ha7 == addr[7:0] ? 8'h0 : _GEN_1266; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1268 = 8'ha8 == addr[7:0] ? 8'h0 : _GEN_1267; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1269 = 8'ha9 == addr[7:0] ? 8'h0 : _GEN_1268; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1270 = 8'haa == addr[7:0] ? 8'h0 : _GEN_1269; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1271 = 8'hab == addr[7:0] ? 8'h0 : _GEN_1270; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1272 = 8'hac == addr[7:0] ? 8'h0 : _GEN_1271; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1273 = 8'had == addr[7:0] ? 8'h0 : _GEN_1272; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1274 = 8'hae == addr[7:0] ? 8'h0 : _GEN_1273; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1275 = 8'haf == addr[7:0] ? 8'h0 : _GEN_1274; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1276 = 8'hb0 == addr[7:0] ? 8'h0 : _GEN_1275; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1277 = 8'hb1 == addr[7:0] ? 8'h0 : _GEN_1276; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1278 = 8'hb2 == addr[7:0] ? 8'h0 : _GEN_1277; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1279 = 8'hb3 == addr[7:0] ? 8'h0 : _GEN_1278; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1280 = 8'hb4 == addr[7:0] ? 8'h0 : _GEN_1279; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1281 = 8'hb5 == addr[7:0] ? 8'h0 : _GEN_1280; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1282 = 8'hb6 == addr[7:0] ? 8'h0 : _GEN_1281; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1283 = 8'hb7 == addr[7:0] ? 8'h0 : _GEN_1282; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1284 = 8'hb8 == addr[7:0] ? 8'h0 : _GEN_1283; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1285 = 8'hb9 == addr[7:0] ? 8'h0 : _GEN_1284; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1286 = 8'hba == addr[7:0] ? 8'h0 : _GEN_1285; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1287 = 8'hbb == addr[7:0] ? 8'h0 : _GEN_1286; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1288 = 8'hbc == addr[7:0] ? 8'h0 : _GEN_1287; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1289 = 8'hbd == addr[7:0] ? 8'h0 : _GEN_1288; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1290 = 8'hbe == addr[7:0] ? 8'h0 : _GEN_1289; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1291 = 8'hbf == addr[7:0] ? 8'h0 : _GEN_1290; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1292 = 8'hc0 == addr[7:0] ? 8'h0 : _GEN_1291; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1293 = 8'hc1 == addr[7:0] ? 8'h0 : _GEN_1292; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1294 = 8'hc2 == addr[7:0] ? 8'h0 : _GEN_1293; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1295 = 8'hc3 == addr[7:0] ? 8'h0 : _GEN_1294; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1296 = 8'hc4 == addr[7:0] ? 8'h0 : _GEN_1295; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1297 = 8'hc5 == addr[7:0] ? 8'h0 : _GEN_1296; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1298 = 8'hc6 == addr[7:0] ? 8'h0 : _GEN_1297; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1299 = 8'hc7 == addr[7:0] ? 8'h0 : _GEN_1298; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1300 = 8'hc8 == addr[7:0] ? 8'h0 : _GEN_1299; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1301 = 8'hc9 == addr[7:0] ? 8'h0 : _GEN_1300; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1302 = 8'hca == addr[7:0] ? 8'h0 : _GEN_1301; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1303 = 8'hcb == addr[7:0] ? 8'h0 : _GEN_1302; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1304 = 8'hcc == addr[7:0] ? 8'h0 : _GEN_1303; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1305 = 8'hcd == addr[7:0] ? 8'h0 : _GEN_1304; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1306 = 8'hce == addr[7:0] ? 8'h0 : _GEN_1305; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1307 = 8'hcf == addr[7:0] ? 8'h0 : _GEN_1306; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1308 = 8'hd0 == addr[7:0] ? 8'h0 : _GEN_1307; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1309 = 8'hd1 == addr[7:0] ? 8'h0 : _GEN_1308; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1310 = 8'hd2 == addr[7:0] ? 8'h0 : _GEN_1309; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1311 = 8'hd3 == addr[7:0] ? 8'h0 : _GEN_1310; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1312 = 8'hd4 == addr[7:0] ? 8'h0 : _GEN_1311; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1313 = 8'hd5 == addr[7:0] ? 8'h0 : _GEN_1312; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1314 = 8'hd6 == addr[7:0] ? 8'h0 : _GEN_1313; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1315 = 8'hd7 == addr[7:0] ? 8'h0 : _GEN_1314; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1316 = 8'hd8 == addr[7:0] ? 8'h0 : _GEN_1315; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1317 = 8'hd9 == addr[7:0] ? 8'h0 : _GEN_1316; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1318 = 8'hda == addr[7:0] ? 8'h0 : _GEN_1317; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1319 = 8'hdb == addr[7:0] ? 8'h0 : _GEN_1318; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1321 = 8'h1 == _T_16[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1322 = 8'h2 == _T_16[7:0] ? 8'h0 : _GEN_1321; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1323 = 8'h3 == _T_16[7:0] ? 8'hfe : _GEN_1322; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1324 = 8'h4 == _T_16[7:0] ? 8'h93 : _GEN_1323; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1325 = 8'h5 == _T_16[7:0] ? 8'h5 : _GEN_1324; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1326 = 8'h6 == _T_16[7:0] ? 8'h0 : _GEN_1325; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1327 = 8'h7 == _T_16[7:0] ? 8'hfc : _GEN_1326; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1328 = 8'h8 == _T_16[7:0] ? 8'h33 : _GEN_1327; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1329 = 8'h9 == _T_16[7:0] ? 8'h6 : _GEN_1328; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1330 = 8'ha == _T_16[7:0] ? 8'hb5 : _GEN_1329; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1331 = 8'hb == _T_16[7:0] ? 8'h0 : _GEN_1330; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1332 = 8'hc == _T_16[7:0] ? 8'h13 : _GEN_1331; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1333 = 8'hd == _T_16[7:0] ? 8'h5 : _GEN_1332; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1334 = 8'he == _T_16[7:0] ? 8'ha0 : _GEN_1333; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1335 = 8'hf == _T_16[7:0] ? 8'h0 : _GEN_1334; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1336 = 8'h10 == _T_16[7:0] ? 8'h73 : _GEN_1335; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1337 = 8'h11 == _T_16[7:0] ? 8'h0 : _GEN_1336; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1338 = 8'h12 == _T_16[7:0] ? 8'h0 : _GEN_1337; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1339 = 8'h13 == _T_16[7:0] ? 8'h0 : _GEN_1338; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1340 = 8'h14 == _T_16[7:0] ? 8'h0 : _GEN_1339; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1341 = 8'h15 == _T_16[7:0] ? 8'h0 : _GEN_1340; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1342 = 8'h16 == _T_16[7:0] ? 8'h0 : _GEN_1341; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1343 = 8'h17 == _T_16[7:0] ? 8'h0 : _GEN_1342; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1344 = 8'h18 == _T_16[7:0] ? 8'h0 : _GEN_1343; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1345 = 8'h19 == _T_16[7:0] ? 8'h0 : _GEN_1344; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1346 = 8'h1a == _T_16[7:0] ? 8'h0 : _GEN_1345; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1347 = 8'h1b == _T_16[7:0] ? 8'h0 : _GEN_1346; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1348 = 8'h1c == _T_16[7:0] ? 8'h0 : _GEN_1347; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1349 = 8'h1d == _T_16[7:0] ? 8'h0 : _GEN_1348; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1350 = 8'h1e == _T_16[7:0] ? 8'h0 : _GEN_1349; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1351 = 8'h1f == _T_16[7:0] ? 8'h0 : _GEN_1350; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1352 = 8'h20 == _T_16[7:0] ? 8'h0 : _GEN_1351; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1353 = 8'h21 == _T_16[7:0] ? 8'h0 : _GEN_1352; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1354 = 8'h22 == _T_16[7:0] ? 8'h0 : _GEN_1353; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1355 = 8'h23 == _T_16[7:0] ? 8'h0 : _GEN_1354; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1356 = 8'h24 == _T_16[7:0] ? 8'h0 : _GEN_1355; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1357 = 8'h25 == _T_16[7:0] ? 8'h0 : _GEN_1356; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1358 = 8'h26 == _T_16[7:0] ? 8'h0 : _GEN_1357; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1359 = 8'h27 == _T_16[7:0] ? 8'h0 : _GEN_1358; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1360 = 8'h28 == _T_16[7:0] ? 8'h0 : _GEN_1359; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1361 = 8'h29 == _T_16[7:0] ? 8'h0 : _GEN_1360; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1362 = 8'h2a == _T_16[7:0] ? 8'h0 : _GEN_1361; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1363 = 8'h2b == _T_16[7:0] ? 8'h0 : _GEN_1362; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1364 = 8'h2c == _T_16[7:0] ? 8'h0 : _GEN_1363; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1365 = 8'h2d == _T_16[7:0] ? 8'h0 : _GEN_1364; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1366 = 8'h2e == _T_16[7:0] ? 8'h0 : _GEN_1365; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1367 = 8'h2f == _T_16[7:0] ? 8'h0 : _GEN_1366; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1368 = 8'h30 == _T_16[7:0] ? 8'h0 : _GEN_1367; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1369 = 8'h31 == _T_16[7:0] ? 8'h0 : _GEN_1368; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1370 = 8'h32 == _T_16[7:0] ? 8'h0 : _GEN_1369; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1371 = 8'h33 == _T_16[7:0] ? 8'h0 : _GEN_1370; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1372 = 8'h34 == _T_16[7:0] ? 8'h0 : _GEN_1371; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1373 = 8'h35 == _T_16[7:0] ? 8'h0 : _GEN_1372; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1374 = 8'h36 == _T_16[7:0] ? 8'h0 : _GEN_1373; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1375 = 8'h37 == _T_16[7:0] ? 8'h0 : _GEN_1374; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1376 = 8'h38 == _T_16[7:0] ? 8'h0 : _GEN_1375; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1377 = 8'h39 == _T_16[7:0] ? 8'h0 : _GEN_1376; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1378 = 8'h3a == _T_16[7:0] ? 8'h0 : _GEN_1377; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1379 = 8'h3b == _T_16[7:0] ? 8'h0 : _GEN_1378; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1380 = 8'h3c == _T_16[7:0] ? 8'h0 : _GEN_1379; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1381 = 8'h3d == _T_16[7:0] ? 8'h0 : _GEN_1380; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1382 = 8'h3e == _T_16[7:0] ? 8'h0 : _GEN_1381; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1383 = 8'h3f == _T_16[7:0] ? 8'h0 : _GEN_1382; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1384 = 8'h40 == _T_16[7:0] ? 8'h0 : _GEN_1383; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1385 = 8'h41 == _T_16[7:0] ? 8'h0 : _GEN_1384; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1386 = 8'h42 == _T_16[7:0] ? 8'h0 : _GEN_1385; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1387 = 8'h43 == _T_16[7:0] ? 8'h0 : _GEN_1386; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1388 = 8'h44 == _T_16[7:0] ? 8'h0 : _GEN_1387; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1389 = 8'h45 == _T_16[7:0] ? 8'h0 : _GEN_1388; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1390 = 8'h46 == _T_16[7:0] ? 8'h0 : _GEN_1389; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1391 = 8'h47 == _T_16[7:0] ? 8'h0 : _GEN_1390; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1392 = 8'h48 == _T_16[7:0] ? 8'h0 : _GEN_1391; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1393 = 8'h49 == _T_16[7:0] ? 8'h0 : _GEN_1392; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1394 = 8'h4a == _T_16[7:0] ? 8'h0 : _GEN_1393; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1395 = 8'h4b == _T_16[7:0] ? 8'h0 : _GEN_1394; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1396 = 8'h4c == _T_16[7:0] ? 8'h0 : _GEN_1395; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1397 = 8'h4d == _T_16[7:0] ? 8'h0 : _GEN_1396; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1398 = 8'h4e == _T_16[7:0] ? 8'h0 : _GEN_1397; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1399 = 8'h4f == _T_16[7:0] ? 8'h0 : _GEN_1398; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1400 = 8'h50 == _T_16[7:0] ? 8'h0 : _GEN_1399; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1401 = 8'h51 == _T_16[7:0] ? 8'h0 : _GEN_1400; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1402 = 8'h52 == _T_16[7:0] ? 8'h0 : _GEN_1401; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1403 = 8'h53 == _T_16[7:0] ? 8'h0 : _GEN_1402; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1404 = 8'h54 == _T_16[7:0] ? 8'h0 : _GEN_1403; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1405 = 8'h55 == _T_16[7:0] ? 8'h0 : _GEN_1404; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1406 = 8'h56 == _T_16[7:0] ? 8'h0 : _GEN_1405; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1407 = 8'h57 == _T_16[7:0] ? 8'h0 : _GEN_1406; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1408 = 8'h58 == _T_16[7:0] ? 8'h0 : _GEN_1407; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1409 = 8'h59 == _T_16[7:0] ? 8'h0 : _GEN_1408; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1410 = 8'h5a == _T_16[7:0] ? 8'h0 : _GEN_1409; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1411 = 8'h5b == _T_16[7:0] ? 8'h0 : _GEN_1410; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1412 = 8'h5c == _T_16[7:0] ? 8'h0 : _GEN_1411; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1413 = 8'h5d == _T_16[7:0] ? 8'h0 : _GEN_1412; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1414 = 8'h5e == _T_16[7:0] ? 8'h0 : _GEN_1413; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1415 = 8'h5f == _T_16[7:0] ? 8'h0 : _GEN_1414; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1416 = 8'h60 == _T_16[7:0] ? 8'h0 : _GEN_1415; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1417 = 8'h61 == _T_16[7:0] ? 8'h0 : _GEN_1416; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1418 = 8'h62 == _T_16[7:0] ? 8'h0 : _GEN_1417; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1419 = 8'h63 == _T_16[7:0] ? 8'h0 : _GEN_1418; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1420 = 8'h64 == _T_16[7:0] ? 8'h0 : _GEN_1419; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1421 = 8'h65 == _T_16[7:0] ? 8'h0 : _GEN_1420; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1422 = 8'h66 == _T_16[7:0] ? 8'h0 : _GEN_1421; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1423 = 8'h67 == _T_16[7:0] ? 8'h0 : _GEN_1422; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1424 = 8'h68 == _T_16[7:0] ? 8'h0 : _GEN_1423; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1425 = 8'h69 == _T_16[7:0] ? 8'h0 : _GEN_1424; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1426 = 8'h6a == _T_16[7:0] ? 8'h0 : _GEN_1425; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1427 = 8'h6b == _T_16[7:0] ? 8'h0 : _GEN_1426; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1428 = 8'h6c == _T_16[7:0] ? 8'h0 : _GEN_1427; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1429 = 8'h6d == _T_16[7:0] ? 8'h0 : _GEN_1428; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1430 = 8'h6e == _T_16[7:0] ? 8'h0 : _GEN_1429; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1431 = 8'h6f == _T_16[7:0] ? 8'h0 : _GEN_1430; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1432 = 8'h70 == _T_16[7:0] ? 8'h0 : _GEN_1431; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1433 = 8'h71 == _T_16[7:0] ? 8'h0 : _GEN_1432; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1434 = 8'h72 == _T_16[7:0] ? 8'h0 : _GEN_1433; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1435 = 8'h73 == _T_16[7:0] ? 8'h0 : _GEN_1434; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1436 = 8'h74 == _T_16[7:0] ? 8'h0 : _GEN_1435; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1437 = 8'h75 == _T_16[7:0] ? 8'h0 : _GEN_1436; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1438 = 8'h76 == _T_16[7:0] ? 8'h0 : _GEN_1437; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1439 = 8'h77 == _T_16[7:0] ? 8'h0 : _GEN_1438; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1440 = 8'h78 == _T_16[7:0] ? 8'h0 : _GEN_1439; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1441 = 8'h79 == _T_16[7:0] ? 8'h0 : _GEN_1440; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1442 = 8'h7a == _T_16[7:0] ? 8'h0 : _GEN_1441; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1443 = 8'h7b == _T_16[7:0] ? 8'h0 : _GEN_1442; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1444 = 8'h7c == _T_16[7:0] ? 8'h0 : _GEN_1443; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1445 = 8'h7d == _T_16[7:0] ? 8'h0 : _GEN_1444; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1446 = 8'h7e == _T_16[7:0] ? 8'h0 : _GEN_1445; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1447 = 8'h7f == _T_16[7:0] ? 8'h0 : _GEN_1446; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1448 = 8'h80 == _T_16[7:0] ? 8'h0 : _GEN_1447; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1449 = 8'h81 == _T_16[7:0] ? 8'h0 : _GEN_1448; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1450 = 8'h82 == _T_16[7:0] ? 8'h0 : _GEN_1449; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1451 = 8'h83 == _T_16[7:0] ? 8'h0 : _GEN_1450; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1452 = 8'h84 == _T_16[7:0] ? 8'h0 : _GEN_1451; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1453 = 8'h85 == _T_16[7:0] ? 8'h0 : _GEN_1452; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1454 = 8'h86 == _T_16[7:0] ? 8'h0 : _GEN_1453; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1455 = 8'h87 == _T_16[7:0] ? 8'h0 : _GEN_1454; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1456 = 8'h88 == _T_16[7:0] ? 8'h0 : _GEN_1455; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1457 = 8'h89 == _T_16[7:0] ? 8'h0 : _GEN_1456; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1458 = 8'h8a == _T_16[7:0] ? 8'h0 : _GEN_1457; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1459 = 8'h8b == _T_16[7:0] ? 8'h0 : _GEN_1458; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1460 = 8'h8c == _T_16[7:0] ? 8'h0 : _GEN_1459; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1461 = 8'h8d == _T_16[7:0] ? 8'h0 : _GEN_1460; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1462 = 8'h8e == _T_16[7:0] ? 8'h0 : _GEN_1461; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1463 = 8'h8f == _T_16[7:0] ? 8'h0 : _GEN_1462; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1464 = 8'h90 == _T_16[7:0] ? 8'h0 : _GEN_1463; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1465 = 8'h91 == _T_16[7:0] ? 8'h0 : _GEN_1464; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1466 = 8'h92 == _T_16[7:0] ? 8'h0 : _GEN_1465; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1467 = 8'h93 == _T_16[7:0] ? 8'h0 : _GEN_1466; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1468 = 8'h94 == _T_16[7:0] ? 8'h0 : _GEN_1467; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1469 = 8'h95 == _T_16[7:0] ? 8'h0 : _GEN_1468; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1470 = 8'h96 == _T_16[7:0] ? 8'h0 : _GEN_1469; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1471 = 8'h97 == _T_16[7:0] ? 8'h0 : _GEN_1470; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1472 = 8'h98 == _T_16[7:0] ? 8'h0 : _GEN_1471; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1473 = 8'h99 == _T_16[7:0] ? 8'h0 : _GEN_1472; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1474 = 8'h9a == _T_16[7:0] ? 8'h0 : _GEN_1473; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1475 = 8'h9b == _T_16[7:0] ? 8'h0 : _GEN_1474; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1476 = 8'h9c == _T_16[7:0] ? 8'h0 : _GEN_1475; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1477 = 8'h9d == _T_16[7:0] ? 8'h0 : _GEN_1476; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1478 = 8'h9e == _T_16[7:0] ? 8'h0 : _GEN_1477; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1479 = 8'h9f == _T_16[7:0] ? 8'h0 : _GEN_1478; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1480 = 8'ha0 == _T_16[7:0] ? 8'h0 : _GEN_1479; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1481 = 8'ha1 == _T_16[7:0] ? 8'h0 : _GEN_1480; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1482 = 8'ha2 == _T_16[7:0] ? 8'h0 : _GEN_1481; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1483 = 8'ha3 == _T_16[7:0] ? 8'h0 : _GEN_1482; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1484 = 8'ha4 == _T_16[7:0] ? 8'h0 : _GEN_1483; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1485 = 8'ha5 == _T_16[7:0] ? 8'h0 : _GEN_1484; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1486 = 8'ha6 == _T_16[7:0] ? 8'h0 : _GEN_1485; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1487 = 8'ha7 == _T_16[7:0] ? 8'h0 : _GEN_1486; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1488 = 8'ha8 == _T_16[7:0] ? 8'h0 : _GEN_1487; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1489 = 8'ha9 == _T_16[7:0] ? 8'h0 : _GEN_1488; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1490 = 8'haa == _T_16[7:0] ? 8'h0 : _GEN_1489; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1491 = 8'hab == _T_16[7:0] ? 8'h0 : _GEN_1490; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1492 = 8'hac == _T_16[7:0] ? 8'h0 : _GEN_1491; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1493 = 8'had == _T_16[7:0] ? 8'h0 : _GEN_1492; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1494 = 8'hae == _T_16[7:0] ? 8'h0 : _GEN_1493; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1495 = 8'haf == _T_16[7:0] ? 8'h0 : _GEN_1494; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1496 = 8'hb0 == _T_16[7:0] ? 8'h0 : _GEN_1495; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1497 = 8'hb1 == _T_16[7:0] ? 8'h0 : _GEN_1496; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1498 = 8'hb2 == _T_16[7:0] ? 8'h0 : _GEN_1497; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1499 = 8'hb3 == _T_16[7:0] ? 8'h0 : _GEN_1498; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1500 = 8'hb4 == _T_16[7:0] ? 8'h0 : _GEN_1499; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1501 = 8'hb5 == _T_16[7:0] ? 8'h0 : _GEN_1500; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1502 = 8'hb6 == _T_16[7:0] ? 8'h0 : _GEN_1501; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1503 = 8'hb7 == _T_16[7:0] ? 8'h0 : _GEN_1502; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1504 = 8'hb8 == _T_16[7:0] ? 8'h0 : _GEN_1503; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1505 = 8'hb9 == _T_16[7:0] ? 8'h0 : _GEN_1504; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1506 = 8'hba == _T_16[7:0] ? 8'h0 : _GEN_1505; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1507 = 8'hbb == _T_16[7:0] ? 8'h0 : _GEN_1506; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1508 = 8'hbc == _T_16[7:0] ? 8'h0 : _GEN_1507; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1509 = 8'hbd == _T_16[7:0] ? 8'h0 : _GEN_1508; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1510 = 8'hbe == _T_16[7:0] ? 8'h0 : _GEN_1509; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1511 = 8'hbf == _T_16[7:0] ? 8'h0 : _GEN_1510; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1512 = 8'hc0 == _T_16[7:0] ? 8'h0 : _GEN_1511; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1513 = 8'hc1 == _T_16[7:0] ? 8'h0 : _GEN_1512; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1514 = 8'hc2 == _T_16[7:0] ? 8'h0 : _GEN_1513; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1515 = 8'hc3 == _T_16[7:0] ? 8'h0 : _GEN_1514; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1516 = 8'hc4 == _T_16[7:0] ? 8'h0 : _GEN_1515; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1517 = 8'hc5 == _T_16[7:0] ? 8'h0 : _GEN_1516; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1518 = 8'hc6 == _T_16[7:0] ? 8'h0 : _GEN_1517; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1519 = 8'hc7 == _T_16[7:0] ? 8'h0 : _GEN_1518; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1520 = 8'hc8 == _T_16[7:0] ? 8'h0 : _GEN_1519; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1521 = 8'hc9 == _T_16[7:0] ? 8'h0 : _GEN_1520; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1522 = 8'hca == _T_16[7:0] ? 8'h0 : _GEN_1521; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1523 = 8'hcb == _T_16[7:0] ? 8'h0 : _GEN_1522; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1524 = 8'hcc == _T_16[7:0] ? 8'h0 : _GEN_1523; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1525 = 8'hcd == _T_16[7:0] ? 8'h0 : _GEN_1524; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1526 = 8'hce == _T_16[7:0] ? 8'h0 : _GEN_1525; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1527 = 8'hcf == _T_16[7:0] ? 8'h0 : _GEN_1526; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1528 = 8'hd0 == _T_16[7:0] ? 8'h0 : _GEN_1527; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1529 = 8'hd1 == _T_16[7:0] ? 8'h0 : _GEN_1528; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1530 = 8'hd2 == _T_16[7:0] ? 8'h0 : _GEN_1529; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1531 = 8'hd3 == _T_16[7:0] ? 8'h0 : _GEN_1530; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1532 = 8'hd4 == _T_16[7:0] ? 8'h0 : _GEN_1531; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1533 = 8'hd5 == _T_16[7:0] ? 8'h0 : _GEN_1532; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1534 = 8'hd6 == _T_16[7:0] ? 8'h0 : _GEN_1533; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1535 = 8'hd7 == _T_16[7:0] ? 8'h0 : _GEN_1534; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1536 = 8'hd8 == _T_16[7:0] ? 8'h0 : _GEN_1535; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1537 = 8'hd9 == _T_16[7:0] ? 8'h0 : _GEN_1536; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1538 = 8'hda == _T_16[7:0] ? 8'h0 : _GEN_1537; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1539 = 8'hdb == _T_16[7:0] ? 8'h0 : _GEN_1538; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1541 = 8'h1 == _T_20[7:0] ? 8'h5 : 8'h13; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1542 = 8'h2 == _T_20[7:0] ? 8'h0 : _GEN_1541; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1543 = 8'h3 == _T_20[7:0] ? 8'hfe : _GEN_1542; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1544 = 8'h4 == _T_20[7:0] ? 8'h93 : _GEN_1543; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1545 = 8'h5 == _T_20[7:0] ? 8'h5 : _GEN_1544; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1546 = 8'h6 == _T_20[7:0] ? 8'h0 : _GEN_1545; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1547 = 8'h7 == _T_20[7:0] ? 8'hfc : _GEN_1546; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1548 = 8'h8 == _T_20[7:0] ? 8'h33 : _GEN_1547; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1549 = 8'h9 == _T_20[7:0] ? 8'h6 : _GEN_1548; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1550 = 8'ha == _T_20[7:0] ? 8'hb5 : _GEN_1549; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1551 = 8'hb == _T_20[7:0] ? 8'h0 : _GEN_1550; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1552 = 8'hc == _T_20[7:0] ? 8'h13 : _GEN_1551; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1553 = 8'hd == _T_20[7:0] ? 8'h5 : _GEN_1552; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1554 = 8'he == _T_20[7:0] ? 8'ha0 : _GEN_1553; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1555 = 8'hf == _T_20[7:0] ? 8'h0 : _GEN_1554; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1556 = 8'h10 == _T_20[7:0] ? 8'h73 : _GEN_1555; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1557 = 8'h11 == _T_20[7:0] ? 8'h0 : _GEN_1556; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1558 = 8'h12 == _T_20[7:0] ? 8'h0 : _GEN_1557; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1559 = 8'h13 == _T_20[7:0] ? 8'h0 : _GEN_1558; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1560 = 8'h14 == _T_20[7:0] ? 8'h0 : _GEN_1559; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1561 = 8'h15 == _T_20[7:0] ? 8'h0 : _GEN_1560; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1562 = 8'h16 == _T_20[7:0] ? 8'h0 : _GEN_1561; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1563 = 8'h17 == _T_20[7:0] ? 8'h0 : _GEN_1562; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1564 = 8'h18 == _T_20[7:0] ? 8'h0 : _GEN_1563; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1565 = 8'h19 == _T_20[7:0] ? 8'h0 : _GEN_1564; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1566 = 8'h1a == _T_20[7:0] ? 8'h0 : _GEN_1565; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1567 = 8'h1b == _T_20[7:0] ? 8'h0 : _GEN_1566; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1568 = 8'h1c == _T_20[7:0] ? 8'h0 : _GEN_1567; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1569 = 8'h1d == _T_20[7:0] ? 8'h0 : _GEN_1568; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1570 = 8'h1e == _T_20[7:0] ? 8'h0 : _GEN_1569; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1571 = 8'h1f == _T_20[7:0] ? 8'h0 : _GEN_1570; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1572 = 8'h20 == _T_20[7:0] ? 8'h0 : _GEN_1571; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1573 = 8'h21 == _T_20[7:0] ? 8'h0 : _GEN_1572; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1574 = 8'h22 == _T_20[7:0] ? 8'h0 : _GEN_1573; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1575 = 8'h23 == _T_20[7:0] ? 8'h0 : _GEN_1574; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1576 = 8'h24 == _T_20[7:0] ? 8'h0 : _GEN_1575; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1577 = 8'h25 == _T_20[7:0] ? 8'h0 : _GEN_1576; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1578 = 8'h26 == _T_20[7:0] ? 8'h0 : _GEN_1577; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1579 = 8'h27 == _T_20[7:0] ? 8'h0 : _GEN_1578; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1580 = 8'h28 == _T_20[7:0] ? 8'h0 : _GEN_1579; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1581 = 8'h29 == _T_20[7:0] ? 8'h0 : _GEN_1580; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1582 = 8'h2a == _T_20[7:0] ? 8'h0 : _GEN_1581; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1583 = 8'h2b == _T_20[7:0] ? 8'h0 : _GEN_1582; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1584 = 8'h2c == _T_20[7:0] ? 8'h0 : _GEN_1583; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1585 = 8'h2d == _T_20[7:0] ? 8'h0 : _GEN_1584; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1586 = 8'h2e == _T_20[7:0] ? 8'h0 : _GEN_1585; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1587 = 8'h2f == _T_20[7:0] ? 8'h0 : _GEN_1586; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1588 = 8'h30 == _T_20[7:0] ? 8'h0 : _GEN_1587; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1589 = 8'h31 == _T_20[7:0] ? 8'h0 : _GEN_1588; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1590 = 8'h32 == _T_20[7:0] ? 8'h0 : _GEN_1589; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1591 = 8'h33 == _T_20[7:0] ? 8'h0 : _GEN_1590; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1592 = 8'h34 == _T_20[7:0] ? 8'h0 : _GEN_1591; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1593 = 8'h35 == _T_20[7:0] ? 8'h0 : _GEN_1592; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1594 = 8'h36 == _T_20[7:0] ? 8'h0 : _GEN_1593; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1595 = 8'h37 == _T_20[7:0] ? 8'h0 : _GEN_1594; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1596 = 8'h38 == _T_20[7:0] ? 8'h0 : _GEN_1595; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1597 = 8'h39 == _T_20[7:0] ? 8'h0 : _GEN_1596; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1598 = 8'h3a == _T_20[7:0] ? 8'h0 : _GEN_1597; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1599 = 8'h3b == _T_20[7:0] ? 8'h0 : _GEN_1598; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1600 = 8'h3c == _T_20[7:0] ? 8'h0 : _GEN_1599; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1601 = 8'h3d == _T_20[7:0] ? 8'h0 : _GEN_1600; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1602 = 8'h3e == _T_20[7:0] ? 8'h0 : _GEN_1601; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1603 = 8'h3f == _T_20[7:0] ? 8'h0 : _GEN_1602; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1604 = 8'h40 == _T_20[7:0] ? 8'h0 : _GEN_1603; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1605 = 8'h41 == _T_20[7:0] ? 8'h0 : _GEN_1604; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1606 = 8'h42 == _T_20[7:0] ? 8'h0 : _GEN_1605; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1607 = 8'h43 == _T_20[7:0] ? 8'h0 : _GEN_1606; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1608 = 8'h44 == _T_20[7:0] ? 8'h0 : _GEN_1607; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1609 = 8'h45 == _T_20[7:0] ? 8'h0 : _GEN_1608; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1610 = 8'h46 == _T_20[7:0] ? 8'h0 : _GEN_1609; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1611 = 8'h47 == _T_20[7:0] ? 8'h0 : _GEN_1610; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1612 = 8'h48 == _T_20[7:0] ? 8'h0 : _GEN_1611; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1613 = 8'h49 == _T_20[7:0] ? 8'h0 : _GEN_1612; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1614 = 8'h4a == _T_20[7:0] ? 8'h0 : _GEN_1613; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1615 = 8'h4b == _T_20[7:0] ? 8'h0 : _GEN_1614; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1616 = 8'h4c == _T_20[7:0] ? 8'h0 : _GEN_1615; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1617 = 8'h4d == _T_20[7:0] ? 8'h0 : _GEN_1616; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1618 = 8'h4e == _T_20[7:0] ? 8'h0 : _GEN_1617; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1619 = 8'h4f == _T_20[7:0] ? 8'h0 : _GEN_1618; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1620 = 8'h50 == _T_20[7:0] ? 8'h0 : _GEN_1619; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1621 = 8'h51 == _T_20[7:0] ? 8'h0 : _GEN_1620; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1622 = 8'h52 == _T_20[7:0] ? 8'h0 : _GEN_1621; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1623 = 8'h53 == _T_20[7:0] ? 8'h0 : _GEN_1622; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1624 = 8'h54 == _T_20[7:0] ? 8'h0 : _GEN_1623; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1625 = 8'h55 == _T_20[7:0] ? 8'h0 : _GEN_1624; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1626 = 8'h56 == _T_20[7:0] ? 8'h0 : _GEN_1625; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1627 = 8'h57 == _T_20[7:0] ? 8'h0 : _GEN_1626; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1628 = 8'h58 == _T_20[7:0] ? 8'h0 : _GEN_1627; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1629 = 8'h59 == _T_20[7:0] ? 8'h0 : _GEN_1628; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1630 = 8'h5a == _T_20[7:0] ? 8'h0 : _GEN_1629; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1631 = 8'h5b == _T_20[7:0] ? 8'h0 : _GEN_1630; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1632 = 8'h5c == _T_20[7:0] ? 8'h0 : _GEN_1631; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1633 = 8'h5d == _T_20[7:0] ? 8'h0 : _GEN_1632; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1634 = 8'h5e == _T_20[7:0] ? 8'h0 : _GEN_1633; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1635 = 8'h5f == _T_20[7:0] ? 8'h0 : _GEN_1634; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1636 = 8'h60 == _T_20[7:0] ? 8'h0 : _GEN_1635; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1637 = 8'h61 == _T_20[7:0] ? 8'h0 : _GEN_1636; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1638 = 8'h62 == _T_20[7:0] ? 8'h0 : _GEN_1637; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1639 = 8'h63 == _T_20[7:0] ? 8'h0 : _GEN_1638; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1640 = 8'h64 == _T_20[7:0] ? 8'h0 : _GEN_1639; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1641 = 8'h65 == _T_20[7:0] ? 8'h0 : _GEN_1640; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1642 = 8'h66 == _T_20[7:0] ? 8'h0 : _GEN_1641; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1643 = 8'h67 == _T_20[7:0] ? 8'h0 : _GEN_1642; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1644 = 8'h68 == _T_20[7:0] ? 8'h0 : _GEN_1643; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1645 = 8'h69 == _T_20[7:0] ? 8'h0 : _GEN_1644; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1646 = 8'h6a == _T_20[7:0] ? 8'h0 : _GEN_1645; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1647 = 8'h6b == _T_20[7:0] ? 8'h0 : _GEN_1646; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1648 = 8'h6c == _T_20[7:0] ? 8'h0 : _GEN_1647; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1649 = 8'h6d == _T_20[7:0] ? 8'h0 : _GEN_1648; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1650 = 8'h6e == _T_20[7:0] ? 8'h0 : _GEN_1649; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1651 = 8'h6f == _T_20[7:0] ? 8'h0 : _GEN_1650; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1652 = 8'h70 == _T_20[7:0] ? 8'h0 : _GEN_1651; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1653 = 8'h71 == _T_20[7:0] ? 8'h0 : _GEN_1652; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1654 = 8'h72 == _T_20[7:0] ? 8'h0 : _GEN_1653; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1655 = 8'h73 == _T_20[7:0] ? 8'h0 : _GEN_1654; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1656 = 8'h74 == _T_20[7:0] ? 8'h0 : _GEN_1655; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1657 = 8'h75 == _T_20[7:0] ? 8'h0 : _GEN_1656; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1658 = 8'h76 == _T_20[7:0] ? 8'h0 : _GEN_1657; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1659 = 8'h77 == _T_20[7:0] ? 8'h0 : _GEN_1658; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1660 = 8'h78 == _T_20[7:0] ? 8'h0 : _GEN_1659; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1661 = 8'h79 == _T_20[7:0] ? 8'h0 : _GEN_1660; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1662 = 8'h7a == _T_20[7:0] ? 8'h0 : _GEN_1661; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1663 = 8'h7b == _T_20[7:0] ? 8'h0 : _GEN_1662; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1664 = 8'h7c == _T_20[7:0] ? 8'h0 : _GEN_1663; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1665 = 8'h7d == _T_20[7:0] ? 8'h0 : _GEN_1664; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1666 = 8'h7e == _T_20[7:0] ? 8'h0 : _GEN_1665; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1667 = 8'h7f == _T_20[7:0] ? 8'h0 : _GEN_1666; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1668 = 8'h80 == _T_20[7:0] ? 8'h0 : _GEN_1667; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1669 = 8'h81 == _T_20[7:0] ? 8'h0 : _GEN_1668; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1670 = 8'h82 == _T_20[7:0] ? 8'h0 : _GEN_1669; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1671 = 8'h83 == _T_20[7:0] ? 8'h0 : _GEN_1670; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1672 = 8'h84 == _T_20[7:0] ? 8'h0 : _GEN_1671; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1673 = 8'h85 == _T_20[7:0] ? 8'h0 : _GEN_1672; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1674 = 8'h86 == _T_20[7:0] ? 8'h0 : _GEN_1673; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1675 = 8'h87 == _T_20[7:0] ? 8'h0 : _GEN_1674; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1676 = 8'h88 == _T_20[7:0] ? 8'h0 : _GEN_1675; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1677 = 8'h89 == _T_20[7:0] ? 8'h0 : _GEN_1676; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1678 = 8'h8a == _T_20[7:0] ? 8'h0 : _GEN_1677; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1679 = 8'h8b == _T_20[7:0] ? 8'h0 : _GEN_1678; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1680 = 8'h8c == _T_20[7:0] ? 8'h0 : _GEN_1679; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1681 = 8'h8d == _T_20[7:0] ? 8'h0 : _GEN_1680; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1682 = 8'h8e == _T_20[7:0] ? 8'h0 : _GEN_1681; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1683 = 8'h8f == _T_20[7:0] ? 8'h0 : _GEN_1682; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1684 = 8'h90 == _T_20[7:0] ? 8'h0 : _GEN_1683; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1685 = 8'h91 == _T_20[7:0] ? 8'h0 : _GEN_1684; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1686 = 8'h92 == _T_20[7:0] ? 8'h0 : _GEN_1685; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1687 = 8'h93 == _T_20[7:0] ? 8'h0 : _GEN_1686; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1688 = 8'h94 == _T_20[7:0] ? 8'h0 : _GEN_1687; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1689 = 8'h95 == _T_20[7:0] ? 8'h0 : _GEN_1688; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1690 = 8'h96 == _T_20[7:0] ? 8'h0 : _GEN_1689; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1691 = 8'h97 == _T_20[7:0] ? 8'h0 : _GEN_1690; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1692 = 8'h98 == _T_20[7:0] ? 8'h0 : _GEN_1691; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1693 = 8'h99 == _T_20[7:0] ? 8'h0 : _GEN_1692; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1694 = 8'h9a == _T_20[7:0] ? 8'h0 : _GEN_1693; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1695 = 8'h9b == _T_20[7:0] ? 8'h0 : _GEN_1694; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1696 = 8'h9c == _T_20[7:0] ? 8'h0 : _GEN_1695; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1697 = 8'h9d == _T_20[7:0] ? 8'h0 : _GEN_1696; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1698 = 8'h9e == _T_20[7:0] ? 8'h0 : _GEN_1697; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1699 = 8'h9f == _T_20[7:0] ? 8'h0 : _GEN_1698; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1700 = 8'ha0 == _T_20[7:0] ? 8'h0 : _GEN_1699; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1701 = 8'ha1 == _T_20[7:0] ? 8'h0 : _GEN_1700; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1702 = 8'ha2 == _T_20[7:0] ? 8'h0 : _GEN_1701; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1703 = 8'ha3 == _T_20[7:0] ? 8'h0 : _GEN_1702; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1704 = 8'ha4 == _T_20[7:0] ? 8'h0 : _GEN_1703; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1705 = 8'ha5 == _T_20[7:0] ? 8'h0 : _GEN_1704; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1706 = 8'ha6 == _T_20[7:0] ? 8'h0 : _GEN_1705; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1707 = 8'ha7 == _T_20[7:0] ? 8'h0 : _GEN_1706; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1708 = 8'ha8 == _T_20[7:0] ? 8'h0 : _GEN_1707; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1709 = 8'ha9 == _T_20[7:0] ? 8'h0 : _GEN_1708; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1710 = 8'haa == _T_20[7:0] ? 8'h0 : _GEN_1709; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1711 = 8'hab == _T_20[7:0] ? 8'h0 : _GEN_1710; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1712 = 8'hac == _T_20[7:0] ? 8'h0 : _GEN_1711; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1713 = 8'had == _T_20[7:0] ? 8'h0 : _GEN_1712; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1714 = 8'hae == _T_20[7:0] ? 8'h0 : _GEN_1713; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1715 = 8'haf == _T_20[7:0] ? 8'h0 : _GEN_1714; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1716 = 8'hb0 == _T_20[7:0] ? 8'h0 : _GEN_1715; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1717 = 8'hb1 == _T_20[7:0] ? 8'h0 : _GEN_1716; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1718 = 8'hb2 == _T_20[7:0] ? 8'h0 : _GEN_1717; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1719 = 8'hb3 == _T_20[7:0] ? 8'h0 : _GEN_1718; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1720 = 8'hb4 == _T_20[7:0] ? 8'h0 : _GEN_1719; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1721 = 8'hb5 == _T_20[7:0] ? 8'h0 : _GEN_1720; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1722 = 8'hb6 == _T_20[7:0] ? 8'h0 : _GEN_1721; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1723 = 8'hb7 == _T_20[7:0] ? 8'h0 : _GEN_1722; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1724 = 8'hb8 == _T_20[7:0] ? 8'h0 : _GEN_1723; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1725 = 8'hb9 == _T_20[7:0] ? 8'h0 : _GEN_1724; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1726 = 8'hba == _T_20[7:0] ? 8'h0 : _GEN_1725; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1727 = 8'hbb == _T_20[7:0] ? 8'h0 : _GEN_1726; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1728 = 8'hbc == _T_20[7:0] ? 8'h0 : _GEN_1727; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1729 = 8'hbd == _T_20[7:0] ? 8'h0 : _GEN_1728; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1730 = 8'hbe == _T_20[7:0] ? 8'h0 : _GEN_1729; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1731 = 8'hbf == _T_20[7:0] ? 8'h0 : _GEN_1730; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1732 = 8'hc0 == _T_20[7:0] ? 8'h0 : _GEN_1731; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1733 = 8'hc1 == _T_20[7:0] ? 8'h0 : _GEN_1732; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1734 = 8'hc2 == _T_20[7:0] ? 8'h0 : _GEN_1733; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1735 = 8'hc3 == _T_20[7:0] ? 8'h0 : _GEN_1734; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1736 = 8'hc4 == _T_20[7:0] ? 8'h0 : _GEN_1735; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1737 = 8'hc5 == _T_20[7:0] ? 8'h0 : _GEN_1736; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1738 = 8'hc6 == _T_20[7:0] ? 8'h0 : _GEN_1737; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1739 = 8'hc7 == _T_20[7:0] ? 8'h0 : _GEN_1738; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1740 = 8'hc8 == _T_20[7:0] ? 8'h0 : _GEN_1739; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1741 = 8'hc9 == _T_20[7:0] ? 8'h0 : _GEN_1740; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1742 = 8'hca == _T_20[7:0] ? 8'h0 : _GEN_1741; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1743 = 8'hcb == _T_20[7:0] ? 8'h0 : _GEN_1742; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1744 = 8'hcc == _T_20[7:0] ? 8'h0 : _GEN_1743; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1745 = 8'hcd == _T_20[7:0] ? 8'h0 : _GEN_1744; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1746 = 8'hce == _T_20[7:0] ? 8'h0 : _GEN_1745; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1747 = 8'hcf == _T_20[7:0] ? 8'h0 : _GEN_1746; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1748 = 8'hd0 == _T_20[7:0] ? 8'h0 : _GEN_1747; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1749 = 8'hd1 == _T_20[7:0] ? 8'h0 : _GEN_1748; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1750 = 8'hd2 == _T_20[7:0] ? 8'h0 : _GEN_1749; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1751 = 8'hd3 == _T_20[7:0] ? 8'h0 : _GEN_1750; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1752 = 8'hd4 == _T_20[7:0] ? 8'h0 : _GEN_1751; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1753 = 8'hd5 == _T_20[7:0] ? 8'h0 : _GEN_1752; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1754 = 8'hd6 == _T_20[7:0] ? 8'h0 : _GEN_1753; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1755 = 8'hd7 == _T_20[7:0] ? 8'h0 : _GEN_1754; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1756 = 8'hd8 == _T_20[7:0] ? 8'h0 : _GEN_1755; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1757 = 8'hd9 == _T_20[7:0] ? 8'h0 : _GEN_1756; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1758 = 8'hda == _T_20[7:0] ? 8'h0 : _GEN_1757; // @[Cat.scala 29:58]
  wire [7:0] _GEN_1759 = 8'hdb == _T_20[7:0] ? 8'h0 : _GEN_1758; // @[Cat.scala 29:58]
  wire [31:0] _T_31 = {_GEN_1539,_GEN_1759,_GEN_1099,_GEN_1319}; // @[Cat.scala 29:58]
  assign sysBusIO_s_rdData = _T_14 ? _T_31 : 32'h0; // @[ROM.scala 27:21 ROM.scala 29:23]
  assign instrBus_instr = {_T_11,_T_10}; // @[ROM.scala 24:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    addr <= sysBusIO_m_addr;
    _T_14 <= sysBusIO_m_cmd == 2'h1;
  end
endmodule
module RAM(
  input         clock,
  input  [1:0]  sysBusIO_m_cmd,
  input  [31:0] sysBusIO_m_addr,
  input  [31:0] sysBusIO_m_wrData,
  input         sysBusIO_m_strb_0,
  input         sysBusIO_m_strb_1,
  input         sysBusIO_m_strb_2,
  input         sysBusIO_m_strb_3,
  output [31:0] sysBusIO_s_rdData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] banks_0 [0:1023]; // @[RAM.scala 9:38]
  wire [7:0] banks_0__T_9_data; // @[RAM.scala 9:38]
  wire [9:0] banks_0__T_9_addr; // @[RAM.scala 9:38]
  wire [7:0] banks_0__T_104_data; // @[RAM.scala 9:38]
  wire [9:0] banks_0__T_104_addr; // @[RAM.scala 9:38]
  wire  banks_0__T_104_mask; // @[RAM.scala 9:38]
  wire  banks_0__T_104_en; // @[RAM.scala 9:38]
  reg [9:0] banks_0__T_9_addr_pipe_0;
  reg [7:0] banks_1 [0:1023]; // @[RAM.scala 9:38]
  wire [7:0] banks_1__T_18_data; // @[RAM.scala 9:38]
  wire [9:0] banks_1__T_18_addr; // @[RAM.scala 9:38]
  wire [7:0] banks_1__T_106_data; // @[RAM.scala 9:38]
  wire [9:0] banks_1__T_106_addr; // @[RAM.scala 9:38]
  wire  banks_1__T_106_mask; // @[RAM.scala 9:38]
  wire  banks_1__T_106_en; // @[RAM.scala 9:38]
  reg [9:0] banks_1__T_18_addr_pipe_0;
  reg [7:0] banks_2 [0:1023]; // @[RAM.scala 9:38]
  wire [7:0] banks_2__T_27_data; // @[RAM.scala 9:38]
  wire [9:0] banks_2__T_27_addr; // @[RAM.scala 9:38]
  wire [7:0] banks_2__T_108_data; // @[RAM.scala 9:38]
  wire [9:0] banks_2__T_108_addr; // @[RAM.scala 9:38]
  wire  banks_2__T_108_mask; // @[RAM.scala 9:38]
  wire  banks_2__T_108_en; // @[RAM.scala 9:38]
  reg [9:0] banks_2__T_27_addr_pipe_0;
  reg [7:0] banks_3 [0:1023]; // @[RAM.scala 9:38]
  wire [7:0] banks_3__T_36_data; // @[RAM.scala 9:38]
  wire [9:0] banks_3__T_36_addr; // @[RAM.scala 9:38]
  wire [7:0] banks_3__T_110_data; // @[RAM.scala 9:38]
  wire [9:0] banks_3__T_110_addr; // @[RAM.scala 9:38]
  wire  banks_3__T_110_mask; // @[RAM.scala 9:38]
  wire  banks_3__T_110_en; // @[RAM.scala 9:38]
  reg [9:0] banks_3__T_36_addr_pipe_0;
  wire [1:0] byteOffset = sysBusIO_m_addr[1:0]; // @[RAM.scala 14:21]
  wire  _T_2 = byteOffset > 2'h0; // @[RAM.scala 16:75]
  wire [29:0] _T_5 = sysBusIO_m_addr[31:2] + 30'h1; // @[RAM.scala 16:94]
  wire [29:0] _T_7 = _T_2 ? _T_5 : sysBusIO_m_addr[31:2]; // @[RAM.scala 16:63]
  wire  _T_11 = byteOffset > 2'h1; // @[RAM.scala 16:75]
  wire [29:0] _T_16 = _T_11 ? _T_5 : sysBusIO_m_addr[31:2]; // @[RAM.scala 16:63]
  wire  _T_20 = byteOffset > 2'h2; // @[RAM.scala 16:75]
  wire [29:0] _T_25 = _T_20 ? _T_5 : sysBusIO_m_addr[31:2]; // @[RAM.scala 16:63]
  reg  _T_38; // @[RAM.scala 19:15]
  wire [2:0] _T_39 = {{1'd0}, byteOffset}; // @[RAM.scala 21:88]
  wire [1:0] _T_42 = byteOffset + 2'h1; // @[RAM.scala 21:88]
  wire [1:0] _T_44 = byteOffset + 2'h2; // @[RAM.scala 21:88]
  wire [1:0] _T_46 = byteOffset + 2'h3; // @[RAM.scala 21:88]
  wire [7:0] rdPorts_0 = banks_0__T_9_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] rdPorts_1 = banks_1__T_18_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] _GEN_1 = 2'h1 == _T_39[1:0] ? rdPorts_1 : rdPorts_0; // @[RAM.scala 21:47]
  wire [7:0] rdPorts_2 = banks_2__T_27_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] _GEN_2 = 2'h2 == _T_39[1:0] ? rdPorts_2 : _GEN_1; // @[RAM.scala 21:47]
  wire [7:0] rdPorts_3 = banks_3__T_36_data; // @[RAM.scala 16:24 RAM.scala 16:24]
  wire [7:0] _GEN_3 = 2'h3 == _T_39[1:0] ? rdPorts_3 : _GEN_2; // @[RAM.scala 21:47]
  wire [7:0] _GEN_5 = 2'h1 == _T_42 ? rdPorts_1 : rdPorts_0; // @[RAM.scala 21:47]
  wire [7:0] _GEN_6 = 2'h2 == _T_42 ? rdPorts_2 : _GEN_5; // @[RAM.scala 21:47]
  wire [7:0] _GEN_7 = 2'h3 == _T_42 ? rdPorts_3 : _GEN_6; // @[RAM.scala 21:47]
  wire [7:0] _GEN_9 = 2'h1 == _T_44 ? rdPorts_1 : rdPorts_0; // @[RAM.scala 21:47]
  wire [7:0] _GEN_10 = 2'h2 == _T_44 ? rdPorts_2 : _GEN_9; // @[RAM.scala 21:47]
  wire [7:0] _GEN_11 = 2'h3 == _T_44 ? rdPorts_3 : _GEN_10; // @[RAM.scala 21:47]
  wire [7:0] _GEN_13 = 2'h1 == _T_46 ? rdPorts_1 : rdPorts_0; // @[RAM.scala 21:47]
  wire [7:0] _GEN_14 = 2'h2 == _T_46 ? rdPorts_2 : _GEN_13; // @[RAM.scala 21:47]
  wire [7:0] _GEN_15 = 2'h3 == _T_46 ? rdPorts_3 : _GEN_14; // @[RAM.scala 21:47]
  wire [31:0] _T_50 = {_GEN_15,_GEN_11,_GEN_7,_GEN_3}; // @[Cat.scala 29:58]
  wire [7:0] wrDataInVec_3 = sysBusIO_m_wrData[7:0]; // @[RAM.scala 24:79]
  wire [7:0] wrDataInVec_2 = sysBusIO_m_wrData[15:8]; // @[RAM.scala 24:79]
  wire [7:0] wrDataInVec_1 = sysBusIO_m_wrData[23:16]; // @[RAM.scala 24:79]
  wire [7:0] wrDataInVec_0 = sysBusIO_m_wrData[31:24]; // @[RAM.scala 24:79]
  wire [7:0] _GEN_19 = 2'h1 == _T_46 ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 25:34]
  wire [7:0] _GEN_20 = 2'h2 == _T_46 ? wrDataInVec_2 : _GEN_19; // @[RAM.scala 25:34]
  wire [7:0] _GEN_23 = 2'h1 == _T_44 ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 25:34]
  wire [7:0] _GEN_24 = 2'h2 == _T_44 ? wrDataInVec_2 : _GEN_23; // @[RAM.scala 25:34]
  wire [7:0] _GEN_27 = 2'h1 == _T_42 ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 25:34]
  wire [7:0] _GEN_28 = 2'h2 == _T_42 ? wrDataInVec_2 : _GEN_27; // @[RAM.scala 25:34]
  wire [7:0] _GEN_31 = 2'h1 == _T_39[1:0] ? wrDataInVec_1 : wrDataInVec_0; // @[RAM.scala 25:34]
  wire [7:0] _GEN_32 = 2'h2 == _T_39[1:0] ? wrDataInVec_2 : _GEN_31; // @[RAM.scala 25:34]
  wire  _GEN_35 = 2'h1 == _T_39[1:0] ? sysBusIO_m_strb_1 : sysBusIO_m_strb_0; // @[RAM.scala 26:22]
  wire  _GEN_36 = 2'h2 == _T_39[1:0] ? sysBusIO_m_strb_2 : _GEN_35; // @[RAM.scala 26:22]
  wire  enVec_0 = 2'h3 == _T_39[1:0] ? sysBusIO_m_strb_3 : _GEN_36; // @[RAM.scala 26:22]
  wire  _GEN_39 = 2'h1 == _T_42 ? sysBusIO_m_strb_1 : sysBusIO_m_strb_0; // @[RAM.scala 26:22]
  wire  _GEN_40 = 2'h2 == _T_42 ? sysBusIO_m_strb_2 : _GEN_39; // @[RAM.scala 26:22]
  wire  enVec_1 = 2'h3 == _T_42 ? sysBusIO_m_strb_3 : _GEN_40; // @[RAM.scala 26:22]
  wire  _GEN_43 = 2'h1 == _T_44 ? sysBusIO_m_strb_1 : sysBusIO_m_strb_0; // @[RAM.scala 26:22]
  wire  _GEN_44 = 2'h2 == _T_44 ? sysBusIO_m_strb_2 : _GEN_43; // @[RAM.scala 26:22]
  wire  enVec_2 = 2'h3 == _T_44 ? sysBusIO_m_strb_3 : _GEN_44; // @[RAM.scala 26:22]
  wire  _GEN_47 = 2'h1 == _T_46 ? sysBusIO_m_strb_1 : sysBusIO_m_strb_0; // @[RAM.scala 26:22]
  wire  _GEN_48 = 2'h2 == _T_46 ? sysBusIO_m_strb_2 : _GEN_47; // @[RAM.scala 26:22]
  wire  enVec_3 = 2'h3 == _T_46 ? sysBusIO_m_strb_3 : _GEN_48; // @[RAM.scala 26:22]
  wire  _T_102 = sysBusIO_m_cmd == 2'h2; // @[RAM.scala 31:23]
  assign banks_0__T_9_addr = banks_0__T_9_addr_pipe_0;
  assign banks_0__T_9_data = banks_0[banks_0__T_9_addr]; // @[RAM.scala 9:38]
  assign banks_0__T_104_data = 2'h3 == _T_46 ? wrDataInVec_3 : _GEN_20;
  assign banks_0__T_104_addr = _T_7[9:0];
  assign banks_0__T_104_mask = 1'h1;
  assign banks_0__T_104_en = _T_102 & enVec_0;
  assign banks_1__T_18_addr = banks_1__T_18_addr_pipe_0;
  assign banks_1__T_18_data = banks_1[banks_1__T_18_addr]; // @[RAM.scala 9:38]
  assign banks_1__T_106_data = 2'h3 == _T_44 ? wrDataInVec_3 : _GEN_24;
  assign banks_1__T_106_addr = _T_16[9:0];
  assign banks_1__T_106_mask = 1'h1;
  assign banks_1__T_106_en = _T_102 & enVec_1;
  assign banks_2__T_27_addr = banks_2__T_27_addr_pipe_0;
  assign banks_2__T_27_data = banks_2[banks_2__T_27_addr]; // @[RAM.scala 9:38]
  assign banks_2__T_108_data = 2'h3 == _T_42 ? wrDataInVec_3 : _GEN_28;
  assign banks_2__T_108_addr = _T_25[9:0];
  assign banks_2__T_108_mask = 1'h1;
  assign banks_2__T_108_en = _T_102 & enVec_2;
  assign banks_3__T_36_addr = banks_3__T_36_addr_pipe_0;
  assign banks_3__T_36_data = banks_3[banks_3__T_36_addr]; // @[RAM.scala 9:38]
  assign banks_3__T_110_data = 2'h3 == _T_39[1:0] ? wrDataInVec_3 : _GEN_32;
  assign banks_3__T_110_addr = sysBusIO_m_addr[11:2];
  assign banks_3__T_110_mask = 1'h1;
  assign banks_3__T_110_en = _T_102 & enVec_3;
  assign sysBusIO_s_rdData = _T_38 ? _T_50 : 32'h0; // @[RAM.scala 17:21 RAM.scala 21:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    banks_3[initvar] = _RAND_6[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  banks_0__T_9_addr_pipe_0 = _RAND_1[9:0];
  _RAND_3 = {1{`RANDOM}};
  banks_1__T_18_addr_pipe_0 = _RAND_3[9:0];
  _RAND_5 = {1{`RANDOM}};
  banks_2__T_27_addr_pipe_0 = _RAND_5[9:0];
  _RAND_7 = {1{`RANDOM}};
  banks_3__T_36_addr_pipe_0 = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  _T_38 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(banks_0__T_104_en & banks_0__T_104_mask) begin
      banks_0[banks_0__T_104_addr] <= banks_0__T_104_data; // @[RAM.scala 9:38]
    end
    banks_0__T_9_addr_pipe_0 <= _T_7[9:0];
    if(banks_1__T_106_en & banks_1__T_106_mask) begin
      banks_1[banks_1__T_106_addr] <= banks_1__T_106_data; // @[RAM.scala 9:38]
    end
    banks_1__T_18_addr_pipe_0 <= _T_16[9:0];
    if(banks_2__T_108_en & banks_2__T_108_mask) begin
      banks_2[banks_2__T_108_addr] <= banks_2__T_108_data; // @[RAM.scala 9:38]
    end
    banks_2__T_27_addr_pipe_0 <= _T_25[9:0];
    if(banks_3__T_110_en & banks_3__T_110_mask) begin
      banks_3[banks_3__T_110_addr] <= banks_3__T_110_data; // @[RAM.scala 9:38]
    end
    banks_3__T_36_addr_pipe_0 <= sysBusIO_m_addr[11:2];
    _T_38 <= sysBusIO_m_cmd == 2'h1;
  end
endmodule
module LedVec(
  input         clock,
  input         reset,
  input  [1:0]  sysBusIO_m_cmd,
  input  [31:0] sysBusIO_m_addr,
  input  [31:0] sysBusIO_m_wrData,
  output [31:0] sysBusIO_s_rdData,
  output [15:0] led_led
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] data; // @[LedVec.scala 18:21]
  reg  config_active; // @[LedVec.scala 19:23]
  wire [15:0] _GEN_0 = config_active ? data : 16'h0; // @[LedVec.scala 22:23]
  reg  _T_2; // @[BusModule.scala 68:37]
  reg [31:0] _T_3; // @[BusModule.scala 68:91]
  wire  _T_4 = 32'h2000 == _T_3; // @[Mux.scala 80:60]
  wire [31:0] _T_5 = _T_4 ? {{16'd0}, data} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_6 = 32'h2001 == _T_3; // @[Mux.scala 80:60]
  wire [31:0] _T_7 = _T_6 ? {{31'd0}, config_active} : _T_5; // @[Mux.scala 80:57]
  wire  _T_10 = sysBusIO_m_addr == 32'h0; // @[BusModule.scala 77:40]
  wire  _T_14 = sysBusIO_m_cmd == 2'h2; // @[BusModule.scala 79:58]
  wire  accessors_0_isWritten = _T_10 & _T_14; // @[BusModule.scala 79:40]
  wire  _T_18 = sysBusIO_m_addr == 32'h1; // @[BusModule.scala 77:40]
  wire  accessors_1_isWritten = _T_18 & _T_14; // @[BusModule.scala 79:40]
  wire [15:0] _T_28 = data | 16'h8000; // @[LedVec.scala 34:21]
  assign sysBusIO_s_rdData = _T_2 ? _T_7 : 32'h0; // @[SysBus.scala 70:17 BusModule.scala 68:23]
  assign led_led = accessors_0_isWritten ? _T_28 : _GEN_0; // @[LedVec.scala 23:13 LedVec.scala 25:13 LedVec.scala 34:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  config_active = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      data <= 16'h0;
    end else if (accessors_0_isWritten) begin
      data <= sysBusIO_m_wrData[15:0];
    end
    if (reset) begin
      config_active <= 1'h0;
    end else if (accessors_1_isWritten) begin
      config_active <= sysBusIO_m_wrData[0];
    end
    _T_2 <= sysBusIO_m_cmd == 2'h1;
    _T_3 <= sysBusIO_m_addr;
  end
endmodule
module TypeWriterCore(
  input         clock,
  input         reset,
  output [15:0] led_led
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  pipeline_clock; // @[BareCore.scala 10:24]
  wire  pipeline_reset; // @[BareCore.scala 10:24]
  wire [1:0] pipeline_io_sysBusIO_m_cmd; // @[BareCore.scala 10:24]
  wire [31:0] pipeline_io_sysBusIO_m_addr; // @[BareCore.scala 10:24]
  wire [31:0] pipeline_io_sysBusIO_m_wrData; // @[BareCore.scala 10:24]
  wire  pipeline_io_sysBusIO_m_strb_0; // @[BareCore.scala 10:24]
  wire  pipeline_io_sysBusIO_m_strb_1; // @[BareCore.scala 10:24]
  wire  pipeline_io_sysBusIO_m_strb_2; // @[BareCore.scala 10:24]
  wire  pipeline_io_sysBusIO_m_strb_3; // @[BareCore.scala 10:24]
  wire [31:0] pipeline_io_sysBusIO_s_rdData; // @[BareCore.scala 10:24]
  wire [31:0] pipeline_io_instrBus_pc; // @[BareCore.scala 10:24]
  wire [31:0] pipeline_io_instrBus_instr; // @[BareCore.scala 10:24]
  wire  rom_clock; // @[ROM.scala 11:21]
  wire [1:0] rom_sysBusIO_m_cmd; // @[ROM.scala 11:21]
  wire [31:0] rom_sysBusIO_m_addr; // @[ROM.scala 11:21]
  wire [31:0] rom_sysBusIO_s_rdData; // @[ROM.scala 11:21]
  wire [31:0] rom_instrBus_pc; // @[ROM.scala 11:21]
  wire [31:0] rom_instrBus_instr; // @[ROM.scala 11:21]
  wire  ram_clock; // @[RAM.scala 42:21]
  wire [1:0] ram_sysBusIO_m_cmd; // @[RAM.scala 42:21]
  wire [31:0] ram_sysBusIO_m_addr; // @[RAM.scala 42:21]
  wire [31:0] ram_sysBusIO_m_wrData; // @[RAM.scala 42:21]
  wire  ram_sysBusIO_m_strb_0; // @[RAM.scala 42:21]
  wire  ram_sysBusIO_m_strb_1; // @[RAM.scala 42:21]
  wire  ram_sysBusIO_m_strb_2; // @[RAM.scala 42:21]
  wire  ram_sysBusIO_m_strb_3; // @[RAM.scala 42:21]
  wire [31:0] ram_sysBusIO_s_rdData; // @[RAM.scala 42:21]
  wire  ledm_clock; // @[TypeWriterCore.scala 18:20]
  wire  ledm_reset; // @[TypeWriterCore.scala 18:20]
  wire [1:0] ledm_sysBusIO_m_cmd; // @[TypeWriterCore.scala 18:20]
  wire [31:0] ledm_sysBusIO_m_addr; // @[TypeWriterCore.scala 18:20]
  wire [31:0] ledm_sysBusIO_m_wrData; // @[TypeWriterCore.scala 18:20]
  wire [31:0] ledm_sysBusIO_s_rdData; // @[TypeWriterCore.scala 18:20]
  wire [15:0] ledm_led_led; // @[TypeWriterCore.scala 18:20]
  wire [31:0] sysBus_m_addr = pipeline_io_sysBusIO_m_addr; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire  _T = sysBus_m_addr >= 32'h2000; // @[BusModule.scala 12:44]
  wire  _T_1 = sysBus_m_addr < 32'h2002; // @[BusModule.scala 12:71]
  wire  _T_2 = _T & _T_1; // @[BusModule.scala 12:63]
  wire [1:0] sysBus_m_cmd = pipeline_io_sysBusIO_m_cmd; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire  _T_3 = sysBus_m_cmd != 2'h0; // @[SysBus.scala 27:58]
  wire  _T_4 = _T_2 & _T_3; // @[SysBus.scala 27:44]
  reg  _T_5; // @[SysBus.scala 28:27]
  wire  sysBus_m_strb_0 = pipeline_io_sysBusIO_m_strb_0; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire  sysBus_m_strb_1 = pipeline_io_sysBusIO_m_strb_1; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire  sysBus_m_strb_2 = pipeline_io_sysBusIO_m_strb_2; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire  sysBus_m_strb_3 = pipeline_io_sysBusIO_m_strb_3; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire [31:0] sysBus_m_wrData = pipeline_io_sysBusIO_m_wrData; // @[BareCore.scala 11:20 BareCore.scala 12:10]
  wire [31:0] _GEN_7 = _T_5 ? ledm_sysBusIO_s_rdData : 32'h0; // @[SysBus.scala 33:19]
  wire  _T_6 = sysBus_m_addr >= 32'h1000; // @[BusModule.scala 12:44]
  wire  _T_7 = sysBus_m_addr < 32'h2000; // @[BusModule.scala 12:71]
  wire  _T_8 = _T_6 & _T_7; // @[BusModule.scala 12:63]
  wire  _T_10 = _T_8 & _T_3; // @[SysBus.scala 27:44]
  reg  _T_11; // @[SysBus.scala 28:27]
  wire [31:0] _GEN_16 = _T_11 ? ram_sysBusIO_s_rdData : _GEN_7; // @[SysBus.scala 33:19]
  wire  _T_13 = sysBus_m_addr < 32'hdc; // @[BusModule.scala 12:71]
  wire  _T_16 = _T_13 & _T_3; // @[SysBus.scala 27:44]
  reg  _T_17; // @[SysBus.scala 28:27]
  RVPipeline pipeline ( // @[BareCore.scala 10:24]
    .clock(pipeline_clock),
    .reset(pipeline_reset),
    .io_sysBusIO_m_cmd(pipeline_io_sysBusIO_m_cmd),
    .io_sysBusIO_m_addr(pipeline_io_sysBusIO_m_addr),
    .io_sysBusIO_m_wrData(pipeline_io_sysBusIO_m_wrData),
    .io_sysBusIO_m_strb_0(pipeline_io_sysBusIO_m_strb_0),
    .io_sysBusIO_m_strb_1(pipeline_io_sysBusIO_m_strb_1),
    .io_sysBusIO_m_strb_2(pipeline_io_sysBusIO_m_strb_2),
    .io_sysBusIO_m_strb_3(pipeline_io_sysBusIO_m_strb_3),
    .io_sysBusIO_s_rdData(pipeline_io_sysBusIO_s_rdData),
    .io_instrBus_pc(pipeline_io_instrBus_pc),
    .io_instrBus_instr(pipeline_io_instrBus_instr)
  );
  ROM rom ( // @[ROM.scala 11:21]
    .clock(rom_clock),
    .sysBusIO_m_cmd(rom_sysBusIO_m_cmd),
    .sysBusIO_m_addr(rom_sysBusIO_m_addr),
    .sysBusIO_s_rdData(rom_sysBusIO_s_rdData),
    .instrBus_pc(rom_instrBus_pc),
    .instrBus_instr(rom_instrBus_instr)
  );
  RAM ram ( // @[RAM.scala 42:21]
    .clock(ram_clock),
    .sysBusIO_m_cmd(ram_sysBusIO_m_cmd),
    .sysBusIO_m_addr(ram_sysBusIO_m_addr),
    .sysBusIO_m_wrData(ram_sysBusIO_m_wrData),
    .sysBusIO_m_strb_0(ram_sysBusIO_m_strb_0),
    .sysBusIO_m_strb_1(ram_sysBusIO_m_strb_1),
    .sysBusIO_m_strb_2(ram_sysBusIO_m_strb_2),
    .sysBusIO_m_strb_3(ram_sysBusIO_m_strb_3),
    .sysBusIO_s_rdData(ram_sysBusIO_s_rdData)
  );
  LedVec ledm ( // @[TypeWriterCore.scala 18:20]
    .clock(ledm_clock),
    .reset(ledm_reset),
    .sysBusIO_m_cmd(ledm_sysBusIO_m_cmd),
    .sysBusIO_m_addr(ledm_sysBusIO_m_addr),
    .sysBusIO_m_wrData(ledm_sysBusIO_m_wrData),
    .sysBusIO_s_rdData(ledm_sysBusIO_s_rdData),
    .led_led(ledm_led_led)
  );
  assign led_led = ledm_led_led; // @[TypeWriterCore.scala 19:7]
  assign pipeline_clock = clock;
  assign pipeline_reset = reset;
  assign pipeline_io_sysBusIO_s_rdData = _T_17 ? rom_sysBusIO_s_rdData : _GEN_16; // @[BareCore.scala 12:10]
  assign pipeline_io_instrBus_instr = rom_instrBus_instr; // @[TypeWriterCore.scala 14:24]
  assign rom_clock = clock;
  assign rom_sysBusIO_m_cmd = _T_16 ? sysBus_m_cmd : 2'h0; // @[SysBus.scala 57:14 SysBus.scala 31:23]
  assign rom_sysBusIO_m_addr = _T_16 ? sysBus_m_addr : 32'h0; // @[SysBus.scala 58:15 SysBus.scala 31:23]
  assign rom_instrBus_pc = pipeline_io_instrBus_pc; // @[TypeWriterCore.scala 14:24]
  assign ram_clock = clock;
  assign ram_sysBusIO_m_cmd = _T_10 ? sysBus_m_cmd : 2'h0; // @[SysBus.scala 57:14 SysBus.scala 31:23]
  assign ram_sysBusIO_m_addr = _T_10 ? sysBus_m_addr : 32'h0; // @[SysBus.scala 58:15 SysBus.scala 31:23]
  assign ram_sysBusIO_m_wrData = _T_10 ? sysBus_m_wrData : 32'h0; // @[SysBus.scala 59:17 SysBus.scala 31:23]
  assign ram_sysBusIO_m_strb_0 = _T_10 & sysBus_m_strb_0; // @[SysBus.scala 60:15 SysBus.scala 31:23]
  assign ram_sysBusIO_m_strb_1 = _T_10 & sysBus_m_strb_1; // @[SysBus.scala 60:15 SysBus.scala 31:23]
  assign ram_sysBusIO_m_strb_2 = _T_10 & sysBus_m_strb_2; // @[SysBus.scala 60:15 SysBus.scala 31:23]
  assign ram_sysBusIO_m_strb_3 = _T_10 & sysBus_m_strb_3; // @[SysBus.scala 60:15 SysBus.scala 31:23]
  assign ledm_clock = clock;
  assign ledm_reset = reset;
  assign ledm_sysBusIO_m_cmd = _T_4 ? sysBus_m_cmd : 2'h0; // @[SysBus.scala 57:14 SysBus.scala 31:23]
  assign ledm_sysBusIO_m_addr = _T_4 ? sysBus_m_addr : 32'h0; // @[SysBus.scala 58:15 SysBus.scala 31:23]
  assign ledm_sysBusIO_m_wrData = _T_4 ? sysBus_m_wrData : 32'h0; // @[SysBus.scala 59:17 SysBus.scala 31:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_11 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_17 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_5 <= _T_2 & _T_3;
    _T_11 <= _T_8 & _T_3;
    _T_17 <= _T_13 & _T_3;
  end
endmodule
